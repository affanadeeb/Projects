Five Input AND circuit

.include TSMC_180nm.txt
.option scale=0.09u
.param SUPPLY = 1.8
.param LAMBDA = 0.09u

.param width_P = 8*LAMBDA
.param width_N = 4*LAMBDA

.global gnd vdd

Vdd vdd gnd 'SUPPLY'
vin1 in1 gnd  PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
vin2 in2 gnd  PULSE(0 1.8 0ns 100ps 100ps 40ns 80ns)
vin3 in3 gnd  PULSE(0 1.8 0ns 100ps 100ps 80ns 160ns)
vin4 in4 gnd  PULSE(0 1.8 0ns 100ps 100ps 160ns 320ns)
vin5 in5 gnd  PULSE(0 1.8 0ns 100ps 100ps 320ns 640ns)

M1000 out not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1001 out not_0/in vdd vdd CMOSP w=4 l=2
+  ad=20 pd=18 as=120 ps=108
M1002 not_0/in in1 fiveinputNAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1003 fiveinputNAND_0/a_113_n14# in4 fiveinputNAND_0/a_76_n14# Gnd CMOSN w=4 l=2
+  ad=40 pd=36 as=40 ps=36
M1004 not_0/in in5 vdd fiveinputNAND_0/w_133_0# CMOSP w=4 l=2
+  ad=100 pd=90 as=0 ps=0
M1005 not_0/in in3 vdd fiveinputNAND_0/w_63_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 not_0/in in1 vdd fiveinputNAND_0/w_0_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 gnd in5 fiveinputNAND_0/a_113_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 fiveinputNAND_0/a_76_n14# in3 fiveinputNAND_0/a_45_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1009 fiveinputNAND_0/a_45_n14# in2 fiveinputNAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 vdd in2 not_0/in fiveinputNAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 vdd in4 not_0/in fiveinputNAND_0/w_100_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
C0 vdd vdd 0.05fF
C1 out gnd 0.08fF
C2 fiveinputNAND_0/w_133_0# in5 0.06fF
C3 fiveinputNAND_0/w_32_0# not_0/in 0.03fF
C4 not_0/in gnd 0.01fF
C5 fiveinputNAND_0/a_45_n14# fiveinputNAND_0/a_76_n14# 0.04fF
C6 fiveinputNAND_0/a_6_n14# in1 0.10fF
C7 in2 fiveinputNAND_0/a_45_n14# 0.14fF
C8 out vdd 0.03fF
C9 out vdd 0.13fF
C10 fiveinputNAND_0/a_6_n14# in2 0.04fF
C11 fiveinputNAND_0/a_6_n14# gnd 0.35fF
C12 not_0/in vdd 0.06fF
C13 not_0/in vdd 2.75fF
C14 out not_0/in 0.16fF
C15 vdd fiveinputNAND_0/w_133_0# 0.05fF
C16 fiveinputNAND_0/w_100_0# in4 0.06fF
C17 fiveinputNAND_0/w_100_0# vdd 0.05fF
C18 in1 fiveinputNAND_0/w_0_0# 0.06fF
C19 in3 fiveinputNAND_0/w_63_0# 0.06fF
C20 fiveinputNAND_0/a_6_n14# not_0/in 0.11fF
C21 fiveinputNAND_0/w_63_0# vdd 0.05fF
C22 not_0/in fiveinputNAND_0/w_133_0# 0.03fF
C23 gnd in1 0.20fF
C24 fiveinputNAND_0/a_6_n14# fiveinputNAND_0/a_45_n14# 0.04fF
C25 fiveinputNAND_0/w_32_0# in2 0.06fF
C26 in2 gnd 0.27fF
C27 fiveinputNAND_0/w_100_0# not_0/in 0.03fF
C28 fiveinputNAND_0/a_113_n14# fiveinputNAND_0/a_76_n14# 0.04fF
C29 vdd fiveinputNAND_0/w_0_0# 0.05fF
C30 in3 fiveinputNAND_0/a_76_n14# 0.12fF
C31 fiveinputNAND_0/a_113_n14# gnd 0.04fF
C32 in3 gnd 0.27fF
C33 fiveinputNAND_0/w_63_0# not_0/in 0.03fF
C34 gnd in4 0.26fF
C35 fiveinputNAND_0/a_113_n14# in4 0.14fF
C36 fiveinputNAND_0/w_32_0# vdd 0.05fF
C37 not_0/in fiveinputNAND_0/w_0_0# 0.03fF
C38 out in1 0.04fF
C39 vdd Gnd 0.67fF
C40 fiveinputNAND_0/a_113_n14# Gnd 0.08fF
C41 fiveinputNAND_0/a_76_n14# Gnd 0.05fF
C42 fiveinputNAND_0/a_45_n14# Gnd 0.07fF
C43 fiveinputNAND_0/a_6_n14# Gnd 0.14fF
C44 in5 Gnd 0.15fF
C45 in4 Gnd 0.44fF
C46 in3 Gnd 0.43fF
C47 in2 Gnd 0.39fF
C48 in1 Gnd 0.51fF
C49 fiveinputNAND_0/w_133_0# Gnd 0.43fF
C50 fiveinputNAND_0/w_63_0# Gnd 0.43fF
C51 fiveinputNAND_0/w_32_0# Gnd 0.43fF
C52 fiveinputNAND_0/w_0_0# Gnd 0.43fF
C53 gnd Gnd 0.33fF
C54 out Gnd 0.64fF
C55 not_0/in Gnd 1.48fF
C56 vdd Gnd 0.40fF


.tran 0.1n 800n 
.control
run
set color0 = rgb:f/f/e
set color1 = black
plot v(in1) v(in2)+2 v(in3)+4 v(in4)+6 v(in5)+8 v(out)+10
.end
.endc
