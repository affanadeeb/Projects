magic
tech scmos
timestamp 1699641626
<< nwell >>
rect 0 0 25 16
rect 32 0 57 16
rect 63 0 88 16
<< ntransistor >>
rect 11 -14 13 -10
rect 43 -14 45 -10
rect 74 -14 76 -10
<< ptransistor >>
rect 11 6 13 10
rect 43 6 45 10
rect 74 6 76 10
<< ndiffusion >>
rect 10 -14 11 -10
rect 13 -14 14 -10
rect 42 -14 43 -10
rect 45 -14 46 -10
rect 73 -14 74 -10
rect 76 -14 77 -10
<< pdiffusion >>
rect 10 6 11 10
rect 13 6 14 10
rect 42 6 43 10
rect 45 6 46 10
rect 73 6 74 10
rect 76 6 77 10
<< ndcontact >>
rect 6 -14 10 -10
rect 14 -14 18 -10
rect 38 -14 42 -10
rect 46 -14 50 -10
rect 69 -14 73 -10
rect 77 -14 81 -10
<< pdcontact >>
rect 6 6 10 10
rect 14 6 18 10
rect 38 6 42 10
rect 46 6 50 10
rect 69 6 73 10
rect 77 6 81 10
<< polysilicon >>
rect 11 10 13 13
rect 11 -3 13 6
rect 28 1 30 22
rect 43 10 45 13
rect 74 10 76 13
rect 6 -7 13 -3
rect 11 -10 13 -7
rect 43 -4 45 6
rect 74 -3 76 6
rect 43 -6 49 -4
rect 43 -10 45 -6
rect 74 -7 81 -3
rect 74 -10 76 -7
rect 11 -17 13 -14
rect 43 -17 45 -14
rect 74 -17 76 -14
<< polycontact >>
rect 27 22 31 26
rect 27 -3 31 1
rect 2 -7 6 -3
rect 49 -7 53 -3
rect 81 -7 85 -3
<< metal1 >>
rect 27 26 31 28
rect 31 22 94 25
rect 0 16 88 19
rect 7 10 10 16
rect 46 10 49 16
rect 70 10 73 16
rect 91 10 94 22
rect 81 7 94 10
rect 14 -3 17 6
rect 38 -3 41 6
rect -1 -7 2 -3
rect 14 -6 41 -3
rect 14 -10 17 -6
rect 53 -6 56 -3
rect 85 -7 87 -3
rect 50 -14 69 -11
rect 7 -18 10 -14
rect 38 -18 41 -14
rect 7 -21 41 -18
rect 77 -24 80 -14
rect 0 -27 82 -24
rect 55 -37 60 -35
<< m2contact >>
rect 56 -7 61 -2
rect 55 -35 60 -30
<< metal2 >>
rect 56 -30 59 -7
<< labels >>
rlabel metal1 0 16 57 19 5 vdd
rlabel metal1 0 -7 2 -3 3 in1
rlabel metal1 0 -27 50 -24 1 gnd
rlabel metal1 17 -6 41 -3 1 out
rlabel metal1 85 -7 87 -3 1 in3
rlabel metal1 27 27 31 28 5 out
rlabel metal1 55 -37 60 -35 1 in2
<< end >>
