magic
tech scmos
timestamp 1698585264
<< nwell >>
rect 0 0 25 16
rect 32 0 57 16
<< ntransistor >>
rect 11 -14 13 -10
rect 43 -14 45 -10
<< ptransistor >>
rect 11 6 13 10
rect 43 6 45 10
<< ndiffusion >>
rect 10 -14 11 -10
rect 13 -14 14 -10
rect 42 -14 43 -10
rect 45 -14 46 -10
<< pdiffusion >>
rect 10 6 11 10
rect 13 6 14 10
rect 42 6 43 10
rect 45 6 46 10
<< ndcontact >>
rect 6 -14 10 -10
rect 14 -14 18 -10
rect 38 -14 42 -10
rect 46 -14 50 -10
<< pdcontact >>
rect 6 6 10 10
rect 14 6 18 10
rect 38 6 42 10
rect 46 6 50 10
<< polysilicon >>
rect 11 10 13 13
rect 43 10 45 13
rect 11 -3 13 6
rect 6 -7 13 -3
rect 11 -10 13 -7
rect 43 -4 45 6
rect 43 -6 67 -4
rect 43 -10 45 -6
rect 11 -17 13 -14
rect 43 -17 45 -14
rect 27 -30 30 -19
<< polycontact >>
rect 2 -7 6 -3
rect 67 -7 71 -3
rect 26 -19 31 -14
rect 26 -35 31 -30
<< metal1 >>
rect 0 16 57 19
rect 7 10 10 16
rect 18 6 38 9
rect 50 6 64 9
rect -1 -7 2 -3
rect 18 -14 38 -10
rect 7 -24 10 -14
rect 46 -24 49 -14
rect 7 -27 50 -24
rect 60 -35 64 6
rect 71 -7 74 -3
rect 26 -38 64 -35
<< labels >>
rlabel metal1 0 16 57 19 5 vdd
rlabel metal1 0 -7 2 -3 3 in1
rlabel space 0 -27 50 -24 1 gnd
rlabel metal1 31 -38 60 -35 1 out
rlabel metal1 71 -7 74 -3 7 in2
rlabel metal1 7 -27 49 -24 1 gnd
<< end >>
