magic
tech scmos
timestamp 1699680831
<< metal1 >>
rect 776 261 781 262
rect 867 252 871 254
rect 761 250 820 252
rect 761 249 819 250
rect 621 240 726 243
rect 621 230 624 240
rect 271 227 624 230
rect 638 234 710 237
rect 248 114 262 117
rect 248 106 251 114
rect 271 109 274 227
rect 638 204 641 234
rect 557 201 641 204
rect 261 106 274 109
rect 518 108 547 111
rect 261 84 264 106
rect 557 89 560 201
rect 707 121 710 234
rect 723 129 726 240
rect 761 188 764 249
rect 879 242 882 254
rect 896 229 899 254
rect 982 238 1147 241
rect 982 229 985 238
rect 776 226 818 229
rect 893 226 985 229
rect 998 232 1080 235
rect 776 199 779 226
rect 998 202 1001 232
rect 996 201 1001 202
rect 908 186 944 189
rect 940 175 944 186
rect 1077 176 1080 232
rect 1144 202 1147 238
rect 1144 199 1308 202
rect 1097 187 1143 190
rect 1140 181 1143 187
rect 940 172 983 175
rect 1077 173 1108 176
rect 925 164 974 167
rect 723 126 783 129
rect 707 118 745 121
rect 742 115 745 118
rect 842 115 845 120
rect 742 112 845 115
rect 518 86 560 89
rect 251 81 264 84
rect 885 76 888 121
rect 1105 108 1108 173
rect 1305 161 1308 199
rect 1300 158 1308 161
rect 1137 154 1139 158
rect 1268 127 1341 130
rect 1105 105 1164 108
rect 1161 95 1164 105
rect 885 73 925 76
rect 922 67 925 73
rect 922 64 929 67
rect 451 57 461 60
rect 181 52 192 55
rect 451 51 454 57
rect 744 52 761 55
rect 744 48 747 52
rect 926 35 929 64
rect 1338 53 1341 127
rect 1328 50 1341 53
rect 921 32 929 35
rect 1088 33 1090 36
rect 1111 34 1118 37
rect 188 30 189 32
rect 157 28 160 29
rect 113 25 160 28
rect 181 27 191 30
rect 459 29 462 32
rect 1044 30 1091 33
rect 1131 30 1136 33
rect 389 26 430 29
rect 451 26 462 29
rect 759 26 762 28
rect 683 25 723 26
rect 680 23 723 25
rect 744 23 762 26
rect 1131 22 1134 30
rect 923 17 934 20
rect 1114 19 1135 22
rect 1031 16 1093 19
rect 100 12 160 14
rect 183 12 194 15
rect 376 14 433 15
rect 376 12 430 14
rect 100 11 163 12
rect 5 10 8 11
rect 191 9 199 12
rect 259 9 280 12
rect 453 11 461 14
rect 561 12 571 15
rect 670 11 725 14
rect 722 8 723 11
rect 747 8 761 11
rect 1222 8 1225 16
rect 1252 13 1255 16
rect 1252 10 1311 13
rect 962 5 1225 8
rect 26 -1 31 0
rect 111 -7 114 3
rect 307 1 516 4
rect 303 -18 306 1
rect 601 0 806 3
rect 387 -18 390 -7
rect 596 -27 599 0
rect 803 -3 818 0
rect 850 -9 853 -3
rect 680 -11 685 -9
rect 681 -27 684 -11
rect 752 -26 755 -9
rect 850 -12 947 -9
rect 752 -29 936 -26
rect 933 -31 936 -29
rect 958 -36 961 5
rect 1043 -35 1046 -3
rect 1328 -26 1331 50
rect 1090 -28 1331 -26
rect 1087 -29 1331 -28
rect 1087 -31 1093 -29
<< m2contact >>
rect 776 256 781 261
rect 262 112 268 118
rect 291 113 296 118
rect 547 107 553 113
rect 776 229 781 234
rect 865 201 870 206
rect 996 196 1001 201
rect 1058 175 1063 180
rect 1092 186 1097 191
rect 974 163 979 168
rect 580 109 585 114
rect 927 109 932 114
rect 1132 154 1137 159
rect 1135 132 1140 137
rect 910 57 915 62
rect 429 51 434 56
rect 975 59 982 65
rect 1089 59 1094 64
rect 1118 32 1124 38
rect 110 20 115 25
rect 386 21 391 26
rect 1042 25 1047 30
rect 680 18 685 23
rect 1311 9 1316 14
rect 110 3 115 8
rect 386 -7 391 -2
rect 680 -9 685 -4
rect 751 -9 756 -4
rect 947 -13 952 -8
rect 936 -33 941 -28
rect 1082 -33 1087 -28
<< pm12contact >>
rect 159 52 164 57
<< pdm12contact >>
rect 722 48 727 53
rect 1042 -3 1047 2
<< metal2 >>
rect 777 234 780 256
rect 870 201 931 204
rect 1059 202 1136 205
rect 124 192 127 196
rect 124 189 175 192
rect 172 147 175 189
rect 400 183 403 197
rect 694 186 697 196
rect 694 183 730 186
rect 400 180 435 183
rect 172 144 256 147
rect 253 104 256 144
rect 432 142 435 180
rect 432 139 530 142
rect 268 114 291 117
rect 253 101 273 104
rect 153 54 159 57
rect 269 51 272 101
rect 527 83 530 139
rect 553 109 580 112
rect 527 80 566 83
rect 429 56 432 58
rect 269 48 275 51
rect 111 8 114 20
rect 31 4 38 7
rect 35 -1 38 4
rect 249 -1 252 28
rect 35 -4 252 -1
rect 272 -12 275 48
rect 387 -2 390 21
rect 538 4 545 7
rect 538 -12 541 4
rect 563 -9 566 80
rect 727 69 730 183
rect 928 150 931 201
rect 975 197 996 200
rect 975 168 978 197
rect 1059 187 1092 190
rect 1059 180 1062 187
rect 1044 161 1126 164
rect 928 147 965 150
rect 875 113 878 138
rect 962 134 965 147
rect 1123 136 1126 161
rect 1133 159 1136 202
rect 1123 133 1135 136
rect 1202 127 1210 130
rect 1233 127 1240 130
rect 875 109 927 113
rect 1207 111 1210 127
rect 1237 121 1240 127
rect 1237 118 1345 121
rect 1207 108 1337 111
rect 1091 71 1143 74
rect 727 66 755 69
rect 722 53 725 57
rect 681 -4 684 18
rect 752 -4 755 66
rect 915 59 975 62
rect 1091 64 1094 71
rect 1084 61 1089 64
rect 840 0 849 3
rect 879 0 884 3
rect 1043 2 1046 25
rect 1120 17 1123 32
rect 1334 24 1337 108
rect 1160 20 1167 23
rect 1244 21 1251 24
rect 1160 17 1163 20
rect 1120 14 1163 17
rect 563 -12 642 -9
rect 272 -15 541 -12
rect 538 -20 541 -15
rect 639 -14 642 -12
rect 840 -14 843 0
rect 639 -17 843 -14
rect 538 -21 580 -20
rect 879 -21 882 0
rect 1244 -9 1247 21
rect 952 -12 1247 -9
rect 1282 20 1288 23
rect 1293 21 1337 24
rect 1282 -21 1285 20
rect 1342 13 1345 118
rect 1316 10 1345 13
rect 538 -23 1285 -21
rect 577 -24 1285 -23
rect 941 -32 1082 -29
use XNOR  XNOR_0
timestamp 1699670788
transform 1 0 0 0 1 1
box 0 -1 153 222
use not  not_0
timestamp 1698566035
transform 1 0 159 0 1 33
box 0 -21 25 19
use AND  AND_0
timestamp 1699599481
transform 1 0 193 0 1 8
box -4 1 77 98
use XNOR  XNOR_1
timestamp 1699670788
transform 1 0 276 0 1 2
box 0 -1 153 222
use not  not_1
timestamp 1698566035
transform 1 0 429 0 1 32
box 0 -21 25 19
use threeinputAND  threeinputAND_0
timestamp 1699641646
transform 1 0 460 0 1 2
box -1 -1 101 109
use XNOR  XNOR_2
timestamp 1699670788
transform 1 0 570 0 1 1
box 0 -1 153 222
use not  not_2
timestamp 1698566035
transform 1 0 722 0 1 29
box 0 -21 25 19
use fourinputAND  fourinputAND_0
timestamp 1699642970
transform 1 0 700 0 1 -67
box 59 64 223 130
use fourinputOR  fourinputOR_0
timestamp 1699643964
transform 1 0 785 0 1 123
box -41 -3 140 76
use NOR  NOR_0
timestamp 1698585264
transform 1 0 819 0 1 233
box -1 -38 74 19
use XNOR  XNOR_3
timestamp 1699670788
transform 1 0 931 0 1 6
box 0 -1 153 222
use fourinputAND  fourinputAND_1
timestamp 1699642970
transform 1 0 1079 0 1 59
box 59 64 223 130
use fiveinputAND  fiveinputAND_0
timestamp 1699643694
transform 1 0 1168 0 1 29
box -39 -13 165 67
use not  not_3
timestamp 1698566035
transform 1 0 1089 0 1 40
box 0 -21 25 19
<< labels >>
rlabel metal1 26 -1 31 0 1 A3
rlabel metal1 5 10 8 11 1 gnd
rlabel metal1 111 -7 114 -6 1 B3
rlabel metal1 596 -27 599 -26 1 A1
rlabel metal1 303 -18 306 -17 1 A2
rlabel metal1 387 -18 390 -17 1 B2
rlabel metal1 681 -27 684 -26 1 B1
rlabel metal1 958 -36 961 -35 1 A0
rlabel metal1 1043 -35 1046 -34 1 B0
rlabel metal1 867 252 871 254 5 vdd
rlabel metal1 776 261 781 262 5 greater
rlabel metal1 896 252 899 254 1 Equal
rlabel metal1 879 253 882 254 1 lesser
<< end >>
