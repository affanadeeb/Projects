magic
tech scmos
timestamp 1699782167
<< metal1 >>
rect 947 651 952 652
rect 997 635 1002 636
rect 577 634 582 635
rect 204 618 209 619
rect -166 598 -161 599
rect 1204 577 1270 580
rect 1313 577 1363 580
rect 1204 540 1207 577
rect 1313 555 1348 558
rect 1345 517 1348 555
rect 1360 549 1363 577
rect 1435 562 1440 563
rect 1360 546 1409 549
rect 1237 506 1251 507
rect 1237 504 1252 506
rect 1230 486 1234 487
rect 1230 485 1261 486
rect 1230 484 1262 485
rect 1231 483 1262 484
rect 1321 483 1358 486
rect 2311 453 2314 478
rect 2305 450 2314 453
rect 2131 410 2136 411
rect 2084 385 2157 388
rect 2084 367 2087 385
rect 2227 369 2230 430
rect 2244 369 2247 398
rect 1609 364 2087 367
rect 1609 346 1612 364
rect 2276 362 2279 378
rect 1413 343 1612 346
rect 1314 331 1318 333
rect 1413 331 1416 343
rect 1314 328 1416 331
rect 1314 59 1318 328
rect 2808 206 2811 207
rect 2899 204 2902 205
rect 2993 201 2996 202
rect 3086 198 3089 199
rect 2711 148 2742 150
rect 2711 147 2741 148
rect 1459 107 1462 108
rect 1314 56 1346 59
rect 1474 47 1477 126
rect -198 -198 -195 25
rect -177 -22 -174 22
rect -104 17 -101 22
rect -104 14 -15 17
rect -177 -24 -16 -22
rect -177 -25 -21 -24
rect -3 -58 0 35
rect 16 21 19 46
rect 1412 44 1477 47
rect 189 21 193 22
rect 266 21 269 22
rect 189 19 196 21
rect 12 6 101 9
rect 98 -45 101 6
rect 189 -46 192 19
rect 266 18 290 21
rect 287 -41 290 18
rect 566 11 569 22
rect 383 8 569 11
rect 383 -43 386 8
rect 639 3 642 22
rect 474 0 642 3
rect 474 -43 477 0
rect 936 -9 939 22
rect 564 -12 939 -9
rect 564 -45 567 -12
rect 1009 -24 1012 22
rect 662 -27 1012 -24
rect 1038 -6 1345 -3
rect 662 -51 665 -27
rect 126 -169 134 -166
rect 117 -172 120 -169
rect 131 -183 134 -169
rect 492 -174 495 -167
rect 498 -169 501 -167
rect 498 -172 508 -169
rect 580 -170 583 -164
rect 580 -173 1027 -170
rect -198 -201 1020 -198
rect 109 -226 112 -211
rect 132 -238 135 -212
rect 303 -250 306 -213
rect 320 -262 323 -210
rect 491 -274 494 -209
rect 509 -286 512 -209
rect 1017 -211 1020 -201
rect 1024 -204 1027 -173
rect 1038 -195 1041 -6
rect 1053 -17 1318 -14
rect 1053 -143 1056 -17
rect 1412 -61 1415 44
rect 1491 4 1494 60
rect 1582 33 1585 80
rect 1603 47 1606 98
rect 1651 54 1654 97
rect 1735 61 1738 97
rect 1944 70 1947 88
rect 2029 79 2032 88
rect 2029 76 2242 79
rect 1944 67 2151 70
rect 1735 58 2055 61
rect 1651 51 1957 54
rect 1603 44 1867 47
rect 1582 30 1776 33
rect 1491 1 1724 4
rect 1491 -14 1494 1
rect 1504 -6 1591 -3
rect 1588 -13 1591 -6
rect 1773 -27 1776 30
rect 1864 -27 1867 44
rect 1954 -28 1957 51
rect 2052 -24 2055 58
rect 2148 -25 2151 67
rect 2239 -25 2242 76
rect 2306 78 2309 80
rect 2306 75 2332 78
rect 2329 -26 2332 75
rect 2391 59 2394 80
rect 2391 56 2430 59
rect 2427 -33 2430 56
rect 1608 -42 1729 -39
rect 2711 -41 2714 147
rect 2763 100 2769 104
rect 2819 35 2822 95
rect 2733 32 2822 35
rect 2827 -20 2830 95
rect 2909 91 2912 93
rect 2755 -23 2830 -20
rect 2853 88 2912 91
rect 2920 91 2923 92
rect 2920 88 2952 91
rect 2755 -30 2758 -23
rect 2853 -26 2856 88
rect 2949 -27 2952 88
rect 3004 78 3007 94
rect 3019 90 3022 94
rect 3104 90 3231 93
rect 3019 87 3060 90
rect 3004 75 3043 78
rect 3040 -27 3043 75
rect 3057 65 3060 87
rect 3057 62 3133 65
rect 3130 -28 3133 62
rect 3228 -34 3231 90
rect 1401 -64 1415 -61
rect 1223 -79 1245 -76
rect 1223 -137 1226 -79
rect 3233 -81 3234 -77
rect 1168 -140 1226 -137
rect 1053 -146 1061 -143
rect 1325 -158 1328 -117
rect 1167 -162 1184 -159
rect 1038 -197 1135 -195
rect 1038 -198 1138 -197
rect 1181 -204 1184 -162
rect 1706 -140 1710 -137
rect 1024 -207 1184 -204
rect 1333 -211 1336 -192
rect 678 -298 681 -211
rect 1017 -214 1336 -211
rect 1333 -313 1336 -214
rect 1478 -311 1481 -192
rect 1706 -286 1709 -140
rect 1882 -298 1885 -151
rect 1888 -262 1891 -150
rect 2068 -274 2071 -157
rect 2085 -238 2088 -157
rect 2257 -250 2260 -149
rect 2263 -214 2266 -149
rect 2443 -226 2446 -141
rect 2511 -286 2514 -142
rect 2683 -298 2686 -153
rect 2689 -262 2692 -153
rect 2869 -274 2872 -159
rect 2886 -238 2889 -159
rect 3058 -250 3061 -151
rect 3064 -214 3067 -150
rect 3244 -230 3247 -143
rect 3229 -233 3247 -230
<< m2contact >>
rect 1344 511 1349 517
rect 2131 405 2136 410
rect 1466 400 1471 405
rect 2152 380 2157 385
rect 2141 367 2146 372
rect 2242 421 2247 426
rect 2275 357 2280 362
rect 1394 169 1399 174
rect 1458 102 1463 107
rect 1346 54 1352 60
rect 1602 98 1607 103
rect 1581 80 1586 85
rect 1486 55 1491 60
rect -4 35 1 40
rect -20 9 -15 14
rect -21 -29 -16 -24
rect 15 16 20 21
rect 7 5 12 10
rect 15 -99 20 -94
rect 652 -107 657 -102
rect 667 -153 672 -148
rect -56 -163 -51 -158
rect 677 -164 682 -159
rect 116 -177 121 -172
rect 508 -173 513 -168
rect 302 -180 307 -175
rect 319 -180 324 -175
rect 490 -179 495 -174
rect 131 -188 136 -183
rect 108 -211 113 -206
rect 131 -212 136 -207
rect 108 -231 113 -226
rect 302 -213 307 -208
rect 319 -210 324 -205
rect 490 -209 495 -204
rect 508 -209 513 -204
rect 131 -243 136 -238
rect 303 -255 308 -250
rect 319 -267 324 -262
rect 490 -279 495 -274
rect 677 -211 682 -206
rect 1345 -7 1350 -2
rect 1321 -19 1326 -14
rect 1399 -54 1404 -49
rect 1724 0 1729 5
rect 1499 -7 1504 -2
rect 2737 94 2742 99
rect 2728 31 2733 36
rect 1064 -121 1069 -116
rect 2762 -82 2767 -77
rect 2417 -89 2422 -84
rect 2514 -92 2519 -87
rect 1324 -117 1329 -112
rect 1252 -127 1257 -122
rect 1179 -159 1184 -154
rect 1582 -122 1588 -116
rect 1066 -167 1071 -162
rect 1168 -178 1173 -173
rect 1323 -163 1328 -158
rect 508 -291 513 -286
rect 678 -303 683 -298
rect 1720 -141 1725 -136
rect 2427 -140 2432 -135
rect 1705 -291 1710 -286
rect 1888 -267 1893 -262
rect 2084 -243 2089 -238
rect 2263 -219 2268 -214
rect 2442 -231 2447 -226
rect 2256 -255 2261 -250
rect 2067 -279 2072 -274
rect 2521 -143 2526 -138
rect 2510 -291 2515 -286
rect 2689 -267 2694 -262
rect 2885 -243 2890 -238
rect 3064 -219 3069 -214
rect 3224 -234 3229 -229
rect 3057 -255 3062 -250
rect 2868 -279 2873 -274
rect 1881 -303 1886 -298
rect 2682 -303 2687 -298
<< pdm12contact >>
rect 2762 95 2767 100
<< metal2 >>
rect 1326 369 1329 502
rect 1345 385 1348 511
rect 2141 423 2242 426
rect 1345 382 1383 385
rect 1180 366 1329 369
rect -3 40 0 87
rect -19 6 7 9
rect -20 -50 -17 -29
rect -20 -53 7 -50
rect 16 -94 19 16
rect 657 -106 1068 -103
rect 1065 -116 1068 -106
rect 672 -152 675 -150
rect 672 -155 1062 -152
rect 1180 -154 1183 366
rect 1467 355 1470 400
rect 2133 375 2136 405
rect 2129 372 2136 375
rect 2141 372 2144 423
rect 2153 374 2156 380
rect 2318 374 2321 397
rect 2153 371 2321 374
rect 1322 352 1470 355
rect 1322 -14 1325 352
rect 2276 319 2279 357
rect 1365 170 1394 173
rect 1365 117 1368 170
rect 1334 114 1368 117
rect 1334 -23 1337 114
rect 1436 88 1439 111
rect 1463 103 1607 106
rect 1436 85 1585 88
rect 1352 56 1486 59
rect 2738 56 2741 94
rect 2578 53 2741 56
rect 1729 2 1734 3
rect 1729 0 1788 2
rect 1731 -1 1788 0
rect 1350 -6 1499 -3
rect 1326 -60 1373 -57
rect 1326 -112 1329 -60
rect 1370 -65 1373 -60
rect 1400 -65 1403 -54
rect 1370 -68 1403 -65
rect 1785 -112 1788 -1
rect 2578 -37 2581 53
rect 2725 -33 2728 36
rect 2669 -36 2728 -33
rect 2763 -77 2766 95
rect 2510 -85 2519 -84
rect 2422 -87 2519 -85
rect 2422 -88 2514 -87
rect 1785 -113 1787 -112
rect 1584 -126 1587 -122
rect 1253 -136 1256 -127
rect 1584 -129 1658 -126
rect 1232 -139 1256 -136
rect -56 -219 -53 -163
rect 1059 -163 1062 -155
rect 109 -181 122 -177
rect 109 -206 112 -181
rect 132 -207 135 -188
rect 303 -208 306 -180
rect 320 -205 323 -180
rect 491 -204 494 -179
rect 509 -204 512 -173
rect 678 -206 681 -164
rect 1059 -166 1066 -163
rect 1232 -173 1235 -139
rect 1655 -145 1658 -129
rect 1721 -145 1724 -141
rect 1655 -148 1724 -145
rect 2428 -147 2431 -140
rect 2522 -147 2525 -143
rect 2428 -150 2525 -147
rect 1173 -176 1235 -173
rect 1324 -195 1327 -163
rect 2671 -195 2674 -149
rect 1324 -198 2674 -195
rect -198 -222 3224 -219
rect -198 -234 3224 -231
rect -198 -246 3224 -243
rect -198 -258 3224 -255
rect -198 -270 3224 -267
rect -198 -282 3224 -279
rect -198 -294 3224 -291
rect -198 -306 3224 -303
use addersubtractor  addersubtractor_0
timestamp 1699637881
transform 1 0 -133 0 1 42
box -113 -21 1370 609
use OR  OR_0
timestamp 1699627711
transform 1 0 1063 0 1 -177
box -2 -20 105 58
use enableblock  enableblock_0
timestamp 1699623212
transform 1 0 -46 0 1 -164
box -9 -11 727 123
use AND  AND_2
timestamp 1699599481
transform 1 0 2248 0 1 377
box -4 1 77 98
use twotofourdecoder  twotofourdecoder_0
timestamp 1699604371
transform 1 0 1437 0 1 -179
box -195 -14 172 166
use enableblock  enableblock_1
timestamp 1699623212
transform 1 0 1719 0 1 -146
box -9 -11 727 123
use enableblock  enableblock_2
timestamp 1699623212
transform 1 0 2520 0 1 -148
box -9 -11 727 123
use comparator  comparator_0
timestamp 1699680831
transform 1 0 1348 0 1 115
box 0 -36 1345 262
use AND  AND_0
timestamp 1699599481
transform 1 0 1255 0 1 482
box -4 1 77 98
use XOR  XOR_0
timestamp 1699628355
transform 1 0 1407 0 1 390
box -50 -10 103 172
use andblock  andblock_0
timestamp 1699624517
transform 1 0 2762 0 1 107
box -24 -17 342 99
<< labels >>
rlabel metal1 -166 598 -161 599 1 adder0
rlabel metal1 204 618 209 619 1 adder1
rlabel metal1 577 634 582 635 1 adder2
rlabel metal1 947 651 952 652 5 adder3
rlabel metal1 2808 206 2811 207 1 and3
rlabel metal1 2899 204 2902 205 1 and2
rlabel metal1 2993 201 2996 202 1 and1
rlabel metal1 3086 198 3089 199 1 and0
rlabel metal1 1435 562 1440 563 1 Carry
rlabel metal1 997 635 1002 636 1 vdd
rlabel metal1 3233 -81 3234 -77 1 gnd
rlabel metal1 2311 476 2314 478 1 equal
rlabel metal1 2131 410 2136 411 1 greater
rlabel metal2 -198 -222 -197 -219 1 A0
rlabel metal2 -198 -234 -197 -231 1 B0
rlabel metal2 -198 -246 -197 -243 1 A1
rlabel metal2 -198 -258 -197 -255 1 B1
rlabel metal2 -198 -270 -197 -267 1 A2
rlabel metal2 -198 -282 -197 -279 1 B2
rlabel metal2 -198 -294 -197 -291 1 A3
rlabel metal2 -198 -306 -197 -303 1 B3
rlabel metal1 1333 -313 1336 -312 1 S0
rlabel metal1 1478 -311 1481 -310 1 S1
rlabel metal1 2227 429 2230 430 1 lesser
<< end >>
