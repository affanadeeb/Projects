magic
tech scmos
timestamp 1699643964
<< metal1 >>
rect -10 74 -5 76
rect -14 63 1 66
rect -41 39 -34 43
rect -41 12 -38 39
rect 139 41 140 45
rect 0 35 3 40
rect -13 23 -10 25
rect -13 20 8 23
rect -41 9 27 12
rect -2 0 3 1
rect 99 -2 104 -1
rect 56 -3 61 -2
<< m2contact >>
rect -10 69 -5 74
rect -13 38 -8 43
rect -2 30 3 35
rect -2 1 3 6
<< metal2 >>
rect -9 43 -6 69
rect -8 40 -6 43
rect -1 6 2 30
use not  not_0
timestamp 1698566035
transform 1 0 -35 0 1 46
box 0 -21 25 19
use fourinputNOR  fourinputNOR_0
timestamp 1699185986
transform 1 0 1 0 1 47
box -1 -49 138 19
<< labels >>
rlabel metal1 56 -3 61 -2 1 in2
rlabel metal1 99 -2 104 -1 1 in3
rlabel metal1 139 41 140 45 7 in4
rlabel metal1 -8 63 1 66 5 vdd
rlabel metal1 0 20 8 23 1 gnd
rlabel metal1 -10 74 -5 76 5 out
rlabel metal1 -2 0 3 1 1 in1
<< end >>
