magic
tech scmos
timestamp 1699621976
<< metal1 >>
rect 6 97 11 99
rect 97 97 102 99
rect 187 96 192 98
rect 6 86 54 89
rect 97 88 147 89
rect 97 86 144 88
rect 187 85 240 88
rect 286 66 289 92
rect 283 63 289 66
rect 25 12 35 15
rect -56 -9 -53 12
rect -19 -10 -16 -8
rect 29 -14 32 12
rect 29 -17 103 -14
rect 116 -21 119 15
rect 122 -21 125 15
rect 206 11 221 14
rect 206 -15 209 11
rect 302 -13 305 14
rect 145 -18 210 -15
rect 204 -20 207 -18
<< m2contact >>
rect 6 92 11 97
rect 97 92 102 97
rect 187 91 192 96
rect 6 62 11 67
rect 97 62 102 67
rect 187 61 192 66
rect 14 -9 19 -4
rect 40 -10 45 -5
rect 105 -9 110 -4
rect 103 -19 108 -14
rect 130 -11 135 -6
rect 195 -11 200 -6
rect 140 -19 145 -14
rect 226 -11 231 -6
<< metal2 >>
rect 7 67 10 92
rect 98 67 101 92
rect 188 66 191 91
rect 19 -9 40 -6
rect 110 -9 130 -6
rect 200 -10 226 -7
rect 108 -18 140 -15
use AND  AND_0
timestamp 1699599481
transform 1 0 -52 0 1 -9
box -4 1 77 98
use AND  AND_1
timestamp 1699599481
transform 1 0 39 0 1 -9
box -4 1 77 98
use AND  AND_2
timestamp 1699599481
transform 1 0 129 0 1 -10
box -4 1 77 98
use AND  AND_3
timestamp 1699599481
transform 1 0 225 0 1 -10
box -4 1 77 98
<< labels >>
rlabel metal1 -56 -9 -53 -7 3 in3
rlabel metal1 -19 -10 -16 -8 1 gnd
rlabel metal1 116 -21 119 -20 1 in2
rlabel metal1 122 -21 125 -20 1 in1
rlabel metal1 25 86 32 89 5 vdd
rlabel metal1 204 -20 207 -18 1 enable
rlabel metal1 302 -13 305 -9 7 in0
rlabel metal1 286 91 289 92 5 out0
rlabel metal1 187 96 192 98 5 out1
rlabel metal1 97 97 102 99 5 out2
rlabel metal1 6 97 11 99 5 out3
<< end >>
