NAND gate

.include TSMC_180nm.txt
.option scale=0.09u
.param SUPPLY = 1.8
.param LAMBDA = 0.09u

.param width_P = 8*LAMBDA
.param width_N = 4*LAMBDA

.global vdd

Vdd vdd gnd 'SUPPLY'
vin1 in1 gnd  PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
vin2 in2 gnd  PULSE(0 1.8 0ns 100ps 100ps 40ns 80ns)

M1000 out in1 a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1001 out in1 vdd vdd CMOSP w=4 l=2
+  ad=40 pd=36 as=40 ps=36
M1002 gnd in2 a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1003 vdd in2 out w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
C0 w_32_0# in2 0.06fF
C1 out vdd 0.03fF
C2 vdd out 0.25fF
C3 vdd vdd 0.05fF
C4 in1 vdd 0.06fF
C5 a_6_n14# gnd 0.57fF
C6 w_32_0# out 0.03fF
C7 vdd w_32_0# 0.05fF
C8 out a_6_n14# 0.12fF

.tran 0.1n 200n
.control
run
set color0 = rgb:f/f/e
set color1 = black
plot v(in1) v(in2)+2 v(out)+4
.end
.endc
