ALU
.include TSMC_180nm.txt
.option scale=0.09u
.param SUPPLY = 1.8
.param LAMBDA = 0.09u

.param width_P = 8*LAMBDA
.param width_N = 4*LAMBDA

.global vdd

Vdd vdd gnd 'SUPPLY'
V_in_A3 A3 gnd PULSE(1.8 0 0ns 100ps 100ps 20ns 40ns)
V_in_A2 A2 gnd PULSE(1.8 0 0ns 100ps 100ps 80ns 160ns)
V_in_A1 A1 gnd PULSE(1.8 0 0ns 100ps 100ps 40ns 800ns)
V_in_A0 A0 gnd PULSE(1.8 0 0ns 100ps 100ps 160ns 320ns)
V_in_B3 B3 gnd PULSE(1.8 0 0ns 100ps 100ps 40ns 80ns)
V_in_B2 B2 gnd PULSE(1.8 0 0ns 100ps 100ps 20ns 40ns)
V_in_B1 B1 gnd PULSE(1.8 0 0ns 100ps 100ps 160ns 320ns)
V_in_B0 B0 gnd PULSE(1.8 0 0ns 100ps 100ps 40ns 80ns)



V_in_S1 S1 gnd 0
V_in_S0 S0 gnd 1.8


M1000 addersubtractor_0/fulladder_0/AND_0/not_0/in addersubtractor_0/XOR_0/out addersubtractor_0/fulladder_0/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1001 addersubtractor_0/fulladder_0/AND_0/not_0/in addersubtractor_0/XOR_0/out vdd vdd CMOSP w=4 l=2
+  ad=40 pd=36 as=6210 ps=5584
M1002 gnd enableblock_0/A_out3 addersubtractor_0/fulladder_0/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=3880 pd=3492 as=0 ps=0
M1003 vdd enableblock_0/A_out3 addersubtractor_0/fulladder_0/AND_0/not_0/in addersubtractor_0/fulladder_0/AND_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 addersubtractor_0/fulladder_0/OR_0/in2 addersubtractor_0/fulladder_0/AND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1005 addersubtractor_0/fulladder_0/OR_0/in2 addersubtractor_0/fulladder_0/AND_0/not_0/in vdd addersubtractor_0/fulladder_0/AND_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1006 addersubtractor_0/fulladder_0/AND_1/not_0/in S0 addersubtractor_0/fulladder_0/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1007 addersubtractor_0/fulladder_0/AND_1/not_0/in S0 vdd addersubtractor_0/fulladder_0/AND_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1008 gnd addersubtractor_0/fulladder_0/XOR_1/in2 addersubtractor_0/fulladder_0/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 vdd addersubtractor_0/fulladder_0/XOR_1/in2 addersubtractor_0/fulladder_0/AND_1/not_0/in addersubtractor_0/fulladder_0/AND_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 addersubtractor_0/fulladder_0/OR_0/in1 addersubtractor_0/fulladder_0/AND_1/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1011 addersubtractor_0/fulladder_0/OR_0/in1 addersubtractor_0/fulladder_0/AND_1/not_0/in vdd addersubtractor_0/fulladder_0/AND_1/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1012 addersubtractor_0/fulladder_0/XOR_0/NAND_2/in1 enableblock_0/A_out3 addersubtractor_0/fulladder_0/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1013 addersubtractor_0/fulladder_0/XOR_0/NAND_2/in1 enableblock_0/A_out3 vdd addersubtractor_0/fulladder_0/XOR_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1014 gnd addersubtractor_0/XOR_0/out addersubtractor_0/fulladder_0/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1015 vdd addersubtractor_0/XOR_0/out addersubtractor_0/fulladder_0/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_0/XOR_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1016 addersubtractor_0/fulladder_0/XOR_0/NAND_3/in1 enableblock_0/A_out3 addersubtractor_0/fulladder_0/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1017 addersubtractor_0/fulladder_0/XOR_0/NAND_3/in1 enableblock_0/A_out3 vdd addersubtractor_0/fulladder_0/XOR_0/NAND_1/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1018 gnd addersubtractor_0/fulladder_0/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_0/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1019 vdd addersubtractor_0/fulladder_0/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_0/XOR_0/NAND_3/in1 addersubtractor_0/fulladder_0/XOR_0/NAND_1/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1020 addersubtractor_0/fulladder_0/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_0/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_0/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1021 addersubtractor_0/fulladder_0/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_0/XOR_0/NAND_2/in1 vdd addersubtractor_0/fulladder_0/XOR_0/NAND_2/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1022 gnd addersubtractor_0/XOR_0/out addersubtractor_0/fulladder_0/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1023 vdd addersubtractor_0/XOR_0/out addersubtractor_0/fulladder_0/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_0/XOR_0/NAND_2/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1024 addersubtractor_0/fulladder_0/XOR_1/in2 addersubtractor_0/fulladder_0/XOR_0/NAND_3/in1 addersubtractor_0/fulladder_0/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1025 addersubtractor_0/fulladder_0/XOR_1/in2 addersubtractor_0/fulladder_0/XOR_0/NAND_3/in1 vdd addersubtractor_0/fulladder_0/XOR_0/NAND_3/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1026 gnd addersubtractor_0/fulladder_0/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_0/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1027 vdd addersubtractor_0/fulladder_0/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_0/XOR_1/in2 addersubtractor_0/fulladder_0/XOR_0/NAND_3/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1028 addersubtractor_0/fulladder_0/C addersubtractor_0/fulladder_0/OR_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1029 addersubtractor_0/fulladder_0/C addersubtractor_0/fulladder_0/OR_0/NOT_0/in vdd addersubtractor_0/fulladder_0/OR_0/NOT_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1030 addersubtractor_0/fulladder_0/OR_0/NOT_0/in addersubtractor_0/fulladder_0/OR_0/in1 gnd Gnd CMOSN w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1031 addersubtractor_0/fulladder_0/OR_0/NOR_0/a_13_6# addersubtractor_0/fulladder_0/OR_0/in1 vdd addersubtractor_0/fulladder_0/OR_0/NOR_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1032 gnd addersubtractor_0/fulladder_0/OR_0/in2 addersubtractor_0/fulladder_0/OR_0/NOT_0/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1033 addersubtractor_0/fulladder_0/OR_0/NOT_0/in addersubtractor_0/fulladder_0/OR_0/in2 addersubtractor_0/fulladder_0/OR_0/NOR_0/a_13_6# addersubtractor_0/fulladder_0/OR_0/NOR_0/w_32_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1034 addersubtractor_0/fulladder_0/XOR_1/NAND_2/in1 S0 addersubtractor_0/fulladder_0/XOR_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1035 addersubtractor_0/fulladder_0/XOR_1/NAND_2/in1 S0 vdd addersubtractor_0/fulladder_0/XOR_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1036 gnd addersubtractor_0/fulladder_0/XOR_1/in2 addersubtractor_0/fulladder_0/XOR_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1037 vdd addersubtractor_0/fulladder_0/XOR_1/in2 addersubtractor_0/fulladder_0/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_0/XOR_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1038 addersubtractor_0/fulladder_0/XOR_1/NAND_3/in1 S0 addersubtractor_0/fulladder_0/XOR_1/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1039 addersubtractor_0/fulladder_0/XOR_1/NAND_3/in1 S0 vdd addersubtractor_0/fulladder_0/XOR_1/NAND_1/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1040 gnd addersubtractor_0/fulladder_0/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_0/XOR_1/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1041 vdd addersubtractor_0/fulladder_0/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_0/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_0/XOR_1/NAND_1/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1042 addersubtractor_0/fulladder_0/XOR_1/NAND_3/in2 addersubtractor_0/fulladder_0/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_0/XOR_1/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1043 addersubtractor_0/fulladder_0/XOR_1/NAND_3/in2 addersubtractor_0/fulladder_0/XOR_1/NAND_2/in1 vdd addersubtractor_0/fulladder_0/XOR_1/NAND_2/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1044 gnd addersubtractor_0/fulladder_0/XOR_1/in2 addersubtractor_0/fulladder_0/XOR_1/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1045 vdd addersubtractor_0/fulladder_0/XOR_1/in2 addersubtractor_0/fulladder_0/XOR_1/NAND_3/in2 addersubtractor_0/fulladder_0/XOR_1/NAND_2/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1046 adder0 addersubtractor_0/fulladder_0/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_0/XOR_1/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1047 adder0 addersubtractor_0/fulladder_0/XOR_1/NAND_3/in1 vdd addersubtractor_0/fulladder_0/XOR_1/NAND_3/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1048 gnd addersubtractor_0/fulladder_0/XOR_1/NAND_3/in2 addersubtractor_0/fulladder_0/XOR_1/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1049 vdd addersubtractor_0/fulladder_0/XOR_1/NAND_3/in2 adder0 addersubtractor_0/fulladder_0/XOR_1/NAND_3/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1050 addersubtractor_0/fulladder_1/AND_0/not_0/in addersubtractor_0/XOR_1/out addersubtractor_0/fulladder_1/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1051 addersubtractor_0/fulladder_1/AND_0/not_0/in addersubtractor_0/XOR_1/out vdd addersubtractor_0/fulladder_1/AND_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1052 gnd enableblock_0/A_out1 addersubtractor_0/fulladder_1/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1053 vdd enableblock_0/A_out1 addersubtractor_0/fulladder_1/AND_0/not_0/in addersubtractor_0/fulladder_1/AND_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1054 addersubtractor_0/fulladder_1/OR_0/in2 addersubtractor_0/fulladder_1/AND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1055 addersubtractor_0/fulladder_1/OR_0/in2 addersubtractor_0/fulladder_1/AND_0/not_0/in vdd addersubtractor_0/fulladder_1/AND_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1056 addersubtractor_0/fulladder_1/AND_1/not_0/in addersubtractor_0/fulladder_0/C addersubtractor_0/fulladder_1/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1057 addersubtractor_0/fulladder_1/AND_1/not_0/in addersubtractor_0/fulladder_0/C vdd addersubtractor_0/fulladder_1/AND_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1058 gnd addersubtractor_0/fulladder_1/XOR_1/in2 addersubtractor_0/fulladder_1/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1059 vdd addersubtractor_0/fulladder_1/XOR_1/in2 addersubtractor_0/fulladder_1/AND_1/not_0/in addersubtractor_0/fulladder_1/AND_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1060 addersubtractor_0/fulladder_1/OR_0/in1 addersubtractor_0/fulladder_1/AND_1/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1061 addersubtractor_0/fulladder_1/OR_0/in1 addersubtractor_0/fulladder_1/AND_1/not_0/in vdd addersubtractor_0/fulladder_1/AND_1/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1062 addersubtractor_0/fulladder_1/XOR_0/NAND_2/in1 enableblock_0/A_out1 addersubtractor_0/fulladder_1/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1063 addersubtractor_0/fulladder_1/XOR_0/NAND_2/in1 enableblock_0/A_out1 vdd addersubtractor_0/fulladder_1/XOR_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1064 gnd addersubtractor_0/XOR_1/out addersubtractor_0/fulladder_1/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1065 vdd addersubtractor_0/XOR_1/out addersubtractor_0/fulladder_1/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_1/XOR_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1066 addersubtractor_0/fulladder_1/XOR_0/NAND_3/in1 enableblock_0/A_out1 addersubtractor_0/fulladder_1/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1067 addersubtractor_0/fulladder_1/XOR_0/NAND_3/in1 enableblock_0/A_out1 vdd addersubtractor_0/fulladder_1/XOR_0/NAND_1/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1068 gnd addersubtractor_0/fulladder_1/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_1/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1069 vdd addersubtractor_0/fulladder_1/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_1/XOR_0/NAND_3/in1 addersubtractor_0/fulladder_1/XOR_0/NAND_1/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1070 addersubtractor_0/fulladder_1/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_1/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_1/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1071 addersubtractor_0/fulladder_1/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_1/XOR_0/NAND_2/in1 vdd addersubtractor_0/fulladder_1/XOR_0/NAND_2/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1072 gnd addersubtractor_0/XOR_1/out addersubtractor_0/fulladder_1/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1073 vdd addersubtractor_0/XOR_1/out addersubtractor_0/fulladder_1/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_1/XOR_0/NAND_2/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1074 addersubtractor_0/fulladder_1/XOR_1/in2 addersubtractor_0/fulladder_1/XOR_0/NAND_3/in1 addersubtractor_0/fulladder_1/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1075 addersubtractor_0/fulladder_1/XOR_1/in2 addersubtractor_0/fulladder_1/XOR_0/NAND_3/in1 vdd addersubtractor_0/fulladder_1/XOR_0/NAND_3/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1076 gnd addersubtractor_0/fulladder_1/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_1/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1077 vdd addersubtractor_0/fulladder_1/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_1/XOR_1/in2 addersubtractor_0/fulladder_1/XOR_0/NAND_3/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1078 addersubtractor_0/fulladder_1/C addersubtractor_0/fulladder_1/OR_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1079 addersubtractor_0/fulladder_1/C addersubtractor_0/fulladder_1/OR_0/NOT_0/in vdd addersubtractor_0/fulladder_1/OR_0/NOT_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1080 addersubtractor_0/fulladder_1/OR_0/NOT_0/in addersubtractor_0/fulladder_1/OR_0/in1 gnd Gnd CMOSN w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1081 addersubtractor_0/fulladder_1/OR_0/NOR_0/a_13_6# addersubtractor_0/fulladder_1/OR_0/in1 vdd addersubtractor_0/fulladder_1/OR_0/NOR_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1082 gnd addersubtractor_0/fulladder_1/OR_0/in2 addersubtractor_0/fulladder_1/OR_0/NOT_0/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1083 addersubtractor_0/fulladder_1/OR_0/NOT_0/in addersubtractor_0/fulladder_1/OR_0/in2 addersubtractor_0/fulladder_1/OR_0/NOR_0/a_13_6# addersubtractor_0/fulladder_1/OR_0/NOR_0/w_32_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1084 addersubtractor_0/fulladder_1/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_0/C addersubtractor_0/fulladder_1/XOR_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1085 addersubtractor_0/fulladder_1/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_0/C vdd addersubtractor_0/fulladder_1/XOR_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1086 gnd addersubtractor_0/fulladder_1/XOR_1/in2 addersubtractor_0/fulladder_1/XOR_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1087 vdd addersubtractor_0/fulladder_1/XOR_1/in2 addersubtractor_0/fulladder_1/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_1/XOR_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1088 addersubtractor_0/fulladder_1/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_0/C addersubtractor_0/fulladder_1/XOR_1/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1089 addersubtractor_0/fulladder_1/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_0/C vdd addersubtractor_0/fulladder_1/XOR_1/NAND_1/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1090 gnd addersubtractor_0/fulladder_1/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_1/XOR_1/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1091 vdd addersubtractor_0/fulladder_1/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_1/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_1/XOR_1/NAND_1/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1092 addersubtractor_0/fulladder_1/XOR_1/NAND_3/in2 addersubtractor_0/fulladder_1/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_1/XOR_1/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1093 addersubtractor_0/fulladder_1/XOR_1/NAND_3/in2 addersubtractor_0/fulladder_1/XOR_1/NAND_2/in1 vdd addersubtractor_0/fulladder_1/XOR_1/NAND_2/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1094 gnd addersubtractor_0/fulladder_1/XOR_1/in2 addersubtractor_0/fulladder_1/XOR_1/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1095 vdd addersubtractor_0/fulladder_1/XOR_1/in2 addersubtractor_0/fulladder_1/XOR_1/NAND_3/in2 addersubtractor_0/fulladder_1/XOR_1/NAND_2/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1096 adder1 addersubtractor_0/fulladder_1/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_1/XOR_1/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1097 adder1 addersubtractor_0/fulladder_1/XOR_1/NAND_3/in1 vdd addersubtractor_0/fulladder_1/XOR_1/NAND_3/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1098 gnd addersubtractor_0/fulladder_1/XOR_1/NAND_3/in2 addersubtractor_0/fulladder_1/XOR_1/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1099 vdd addersubtractor_0/fulladder_1/XOR_1/NAND_3/in2 adder1 addersubtractor_0/fulladder_1/XOR_1/NAND_3/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1100 addersubtractor_0/fulladder_2/AND_0/not_0/in addersubtractor_0/XOR_2/out addersubtractor_0/fulladder_2/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1101 addersubtractor_0/fulladder_2/AND_0/not_0/in addersubtractor_0/XOR_2/out vdd addersubtractor_0/fulladder_2/AND_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1102 gnd enableblock_0/B_out3 addersubtractor_0/fulladder_2/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1103 vdd enableblock_0/B_out3 addersubtractor_0/fulladder_2/AND_0/not_0/in addersubtractor_0/fulladder_2/AND_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1104 addersubtractor_0/fulladder_2/OR_0/in2 addersubtractor_0/fulladder_2/AND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1105 addersubtractor_0/fulladder_2/OR_0/in2 addersubtractor_0/fulladder_2/AND_0/not_0/in vdd addersubtractor_0/fulladder_2/AND_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1106 addersubtractor_0/fulladder_2/AND_1/not_0/in addersubtractor_0/fulladder_1/C addersubtractor_0/fulladder_2/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1107 addersubtractor_0/fulladder_2/AND_1/not_0/in addersubtractor_0/fulladder_1/C vdd addersubtractor_0/fulladder_2/AND_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1108 gnd addersubtractor_0/fulladder_2/XOR_1/in2 addersubtractor_0/fulladder_2/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1109 vdd addersubtractor_0/fulladder_2/XOR_1/in2 addersubtractor_0/fulladder_2/AND_1/not_0/in addersubtractor_0/fulladder_2/AND_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1110 addersubtractor_0/fulladder_2/OR_0/in1 addersubtractor_0/fulladder_2/AND_1/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1111 addersubtractor_0/fulladder_2/OR_0/in1 addersubtractor_0/fulladder_2/AND_1/not_0/in vdd addersubtractor_0/fulladder_2/AND_1/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1112 addersubtractor_0/fulladder_2/XOR_0/NAND_2/in1 enableblock_0/B_out3 addersubtractor_0/fulladder_2/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1113 addersubtractor_0/fulladder_2/XOR_0/NAND_2/in1 enableblock_0/B_out3 vdd addersubtractor_0/fulladder_2/XOR_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1114 gnd addersubtractor_0/XOR_2/out addersubtractor_0/fulladder_2/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1115 vdd addersubtractor_0/XOR_2/out addersubtractor_0/fulladder_2/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_2/XOR_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1116 addersubtractor_0/fulladder_2/XOR_0/NAND_3/in1 enableblock_0/B_out3 addersubtractor_0/fulladder_2/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1117 addersubtractor_0/fulladder_2/XOR_0/NAND_3/in1 enableblock_0/B_out3 vdd addersubtractor_0/fulladder_2/XOR_0/NAND_1/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1118 gnd addersubtractor_0/fulladder_2/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_2/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1119 vdd addersubtractor_0/fulladder_2/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_2/XOR_0/NAND_3/in1 addersubtractor_0/fulladder_2/XOR_0/NAND_1/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1120 addersubtractor_0/fulladder_2/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_2/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_2/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1121 addersubtractor_0/fulladder_2/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_2/XOR_0/NAND_2/in1 vdd addersubtractor_0/fulladder_2/XOR_0/NAND_2/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1122 gnd addersubtractor_0/XOR_2/out addersubtractor_0/fulladder_2/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1123 vdd addersubtractor_0/XOR_2/out addersubtractor_0/fulladder_2/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_2/XOR_0/NAND_2/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1124 addersubtractor_0/fulladder_2/XOR_1/in2 addersubtractor_0/fulladder_2/XOR_0/NAND_3/in1 addersubtractor_0/fulladder_2/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1125 addersubtractor_0/fulladder_2/XOR_1/in2 addersubtractor_0/fulladder_2/XOR_0/NAND_3/in1 vdd addersubtractor_0/fulladder_2/XOR_0/NAND_3/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1126 gnd addersubtractor_0/fulladder_2/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_2/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1127 vdd addersubtractor_0/fulladder_2/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_2/XOR_1/in2 addersubtractor_0/fulladder_2/XOR_0/NAND_3/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1128 addersubtractor_0/fulladder_2/C addersubtractor_0/fulladder_2/OR_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1129 addersubtractor_0/fulladder_2/C addersubtractor_0/fulladder_2/OR_0/NOT_0/in vdd addersubtractor_0/fulladder_2/OR_0/NOT_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1130 addersubtractor_0/fulladder_2/OR_0/NOT_0/in addersubtractor_0/fulladder_2/OR_0/in1 gnd Gnd CMOSN w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1131 addersubtractor_0/fulladder_2/OR_0/NOR_0/a_13_6# addersubtractor_0/fulladder_2/OR_0/in1 vdd addersubtractor_0/fulladder_2/OR_0/NOR_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1132 gnd addersubtractor_0/fulladder_2/OR_0/in2 addersubtractor_0/fulladder_2/OR_0/NOT_0/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1133 addersubtractor_0/fulladder_2/OR_0/NOT_0/in addersubtractor_0/fulladder_2/OR_0/in2 addersubtractor_0/fulladder_2/OR_0/NOR_0/a_13_6# addersubtractor_0/fulladder_2/OR_0/NOR_0/w_32_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1134 addersubtractor_0/fulladder_2/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_1/C addersubtractor_0/fulladder_2/XOR_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1135 addersubtractor_0/fulladder_2/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_1/C vdd addersubtractor_0/fulladder_2/XOR_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1136 gnd addersubtractor_0/fulladder_2/XOR_1/in2 addersubtractor_0/fulladder_2/XOR_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1137 vdd addersubtractor_0/fulladder_2/XOR_1/in2 addersubtractor_0/fulladder_2/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_2/XOR_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1138 addersubtractor_0/fulladder_2/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_1/C addersubtractor_0/fulladder_2/XOR_1/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1139 addersubtractor_0/fulladder_2/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_1/C vdd addersubtractor_0/fulladder_2/XOR_1/NAND_1/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1140 gnd addersubtractor_0/fulladder_2/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_2/XOR_1/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1141 vdd addersubtractor_0/fulladder_2/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_2/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_2/XOR_1/NAND_1/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1142 addersubtractor_0/fulladder_2/XOR_1/NAND_3/in2 addersubtractor_0/fulladder_2/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_2/XOR_1/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1143 addersubtractor_0/fulladder_2/XOR_1/NAND_3/in2 addersubtractor_0/fulladder_2/XOR_1/NAND_2/in1 vdd addersubtractor_0/fulladder_2/XOR_1/NAND_2/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1144 gnd addersubtractor_0/fulladder_2/XOR_1/in2 addersubtractor_0/fulladder_2/XOR_1/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1145 vdd addersubtractor_0/fulladder_2/XOR_1/in2 addersubtractor_0/fulladder_2/XOR_1/NAND_3/in2 addersubtractor_0/fulladder_2/XOR_1/NAND_2/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1146 adder2 addersubtractor_0/fulladder_2/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_2/XOR_1/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1147 adder2 addersubtractor_0/fulladder_2/XOR_1/NAND_3/in1 vdd addersubtractor_0/fulladder_2/XOR_1/NAND_3/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1148 gnd addersubtractor_0/fulladder_2/XOR_1/NAND_3/in2 addersubtractor_0/fulladder_2/XOR_1/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1149 vdd addersubtractor_0/fulladder_2/XOR_1/NAND_3/in2 adder2 addersubtractor_0/fulladder_2/XOR_1/NAND_3/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1150 addersubtractor_0/fulladder_3/AND_0/not_0/in addersubtractor_0/XOR_3/out addersubtractor_0/fulladder_3/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1151 addersubtractor_0/fulladder_3/AND_0/not_0/in addersubtractor_0/XOR_3/out vdd addersubtractor_0/fulladder_3/AND_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1152 gnd enableblock_0/B_out1 addersubtractor_0/fulladder_3/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1153 vdd enableblock_0/B_out1 addersubtractor_0/fulladder_3/AND_0/not_0/in addersubtractor_0/fulladder_3/AND_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1154 addersubtractor_0/fulladder_3/OR_0/in2 addersubtractor_0/fulladder_3/AND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1155 addersubtractor_0/fulladder_3/OR_0/in2 addersubtractor_0/fulladder_3/AND_0/not_0/in vdd addersubtractor_0/fulladder_3/AND_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1156 addersubtractor_0/fulladder_3/AND_1/not_0/in addersubtractor_0/fulladder_2/C addersubtractor_0/fulladder_3/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1157 addersubtractor_0/fulladder_3/AND_1/not_0/in addersubtractor_0/fulladder_2/C vdd addersubtractor_0/fulladder_3/AND_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1158 gnd addersubtractor_0/fulladder_3/XOR_1/in2 addersubtractor_0/fulladder_3/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1159 vdd addersubtractor_0/fulladder_3/XOR_1/in2 addersubtractor_0/fulladder_3/AND_1/not_0/in addersubtractor_0/fulladder_3/AND_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1160 addersubtractor_0/fulladder_3/OR_0/in1 addersubtractor_0/fulladder_3/AND_1/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1161 addersubtractor_0/fulladder_3/OR_0/in1 addersubtractor_0/fulladder_3/AND_1/not_0/in vdd addersubtractor_0/fulladder_3/AND_1/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1162 addersubtractor_0/fulladder_3/XOR_0/NAND_2/in1 enableblock_0/B_out1 addersubtractor_0/fulladder_3/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1163 addersubtractor_0/fulladder_3/XOR_0/NAND_2/in1 enableblock_0/B_out1 vdd addersubtractor_0/fulladder_3/XOR_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1164 gnd addersubtractor_0/XOR_3/out addersubtractor_0/fulladder_3/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1165 vdd addersubtractor_0/XOR_3/out addersubtractor_0/fulladder_3/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_3/XOR_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1166 addersubtractor_0/fulladder_3/XOR_0/NAND_3/in1 enableblock_0/B_out1 addersubtractor_0/fulladder_3/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1167 addersubtractor_0/fulladder_3/XOR_0/NAND_3/in1 enableblock_0/B_out1 vdd addersubtractor_0/fulladder_3/XOR_0/NAND_1/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1168 gnd addersubtractor_0/fulladder_3/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_3/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1169 vdd addersubtractor_0/fulladder_3/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_3/XOR_0/NAND_3/in1 addersubtractor_0/fulladder_3/XOR_0/NAND_1/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1170 addersubtractor_0/fulladder_3/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_3/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_3/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1171 addersubtractor_0/fulladder_3/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_3/XOR_0/NAND_2/in1 vdd addersubtractor_0/fulladder_3/XOR_0/NAND_2/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1172 gnd addersubtractor_0/XOR_3/out addersubtractor_0/fulladder_3/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1173 vdd addersubtractor_0/XOR_3/out addersubtractor_0/fulladder_3/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_3/XOR_0/NAND_2/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1174 addersubtractor_0/fulladder_3/XOR_1/in2 addersubtractor_0/fulladder_3/XOR_0/NAND_3/in1 addersubtractor_0/fulladder_3/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1175 addersubtractor_0/fulladder_3/XOR_1/in2 addersubtractor_0/fulladder_3/XOR_0/NAND_3/in1 vdd addersubtractor_0/fulladder_3/XOR_0/NAND_3/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1176 gnd addersubtractor_0/fulladder_3/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_3/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1177 vdd addersubtractor_0/fulladder_3/XOR_0/NAND_3/in2 addersubtractor_0/fulladder_3/XOR_1/in2 addersubtractor_0/fulladder_3/XOR_0/NAND_3/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1178 AND_0/in1 addersubtractor_0/fulladder_3/OR_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1179 AND_0/in1 addersubtractor_0/fulladder_3/OR_0/NOT_0/in vdd addersubtractor_0/fulladder_3/OR_0/NOT_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1180 addersubtractor_0/fulladder_3/OR_0/NOT_0/in addersubtractor_0/fulladder_3/OR_0/in1 gnd Gnd CMOSN w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1181 addersubtractor_0/fulladder_3/OR_0/NOR_0/a_13_6# addersubtractor_0/fulladder_3/OR_0/in1 vdd addersubtractor_0/fulladder_3/OR_0/NOR_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1182 gnd addersubtractor_0/fulladder_3/OR_0/in2 addersubtractor_0/fulladder_3/OR_0/NOT_0/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1183 addersubtractor_0/fulladder_3/OR_0/NOT_0/in addersubtractor_0/fulladder_3/OR_0/in2 addersubtractor_0/fulladder_3/OR_0/NOR_0/a_13_6# addersubtractor_0/fulladder_3/OR_0/NOR_0/w_32_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1184 addersubtractor_0/fulladder_3/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_2/C addersubtractor_0/fulladder_3/XOR_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1185 addersubtractor_0/fulladder_3/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_2/C vdd addersubtractor_0/fulladder_3/XOR_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1186 gnd addersubtractor_0/fulladder_3/XOR_1/in2 addersubtractor_0/fulladder_3/XOR_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1187 vdd addersubtractor_0/fulladder_3/XOR_1/in2 addersubtractor_0/fulladder_3/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_3/XOR_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1188 addersubtractor_0/fulladder_3/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_2/C addersubtractor_0/fulladder_3/XOR_1/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1189 addersubtractor_0/fulladder_3/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_2/C vdd addersubtractor_0/fulladder_3/XOR_1/NAND_1/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1190 gnd addersubtractor_0/fulladder_3/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_3/XOR_1/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1191 vdd addersubtractor_0/fulladder_3/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_3/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_3/XOR_1/NAND_1/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1192 addersubtractor_0/fulladder_3/XOR_1/NAND_3/in2 addersubtractor_0/fulladder_3/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_3/XOR_1/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1193 addersubtractor_0/fulladder_3/XOR_1/NAND_3/in2 addersubtractor_0/fulladder_3/XOR_1/NAND_2/in1 vdd addersubtractor_0/fulladder_3/XOR_1/NAND_2/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1194 gnd addersubtractor_0/fulladder_3/XOR_1/in2 addersubtractor_0/fulladder_3/XOR_1/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1195 vdd addersubtractor_0/fulladder_3/XOR_1/in2 addersubtractor_0/fulladder_3/XOR_1/NAND_3/in2 addersubtractor_0/fulladder_3/XOR_1/NAND_2/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1196 adder3 addersubtractor_0/fulladder_3/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_3/XOR_1/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1197 adder3 addersubtractor_0/fulladder_3/XOR_1/NAND_3/in1 vdd addersubtractor_0/fulladder_3/XOR_1/NAND_3/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1198 gnd addersubtractor_0/fulladder_3/XOR_1/NAND_3/in2 addersubtractor_0/fulladder_3/XOR_1/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1199 vdd addersubtractor_0/fulladder_3/XOR_1/NAND_3/in2 adder3 addersubtractor_0/fulladder_3/XOR_1/NAND_3/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1200 addersubtractor_0/XOR_0/NAND_2/in1 enableblock_0/A_out2 addersubtractor_0/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1201 addersubtractor_0/XOR_0/NAND_2/in1 enableblock_0/A_out2 vdd addersubtractor_0/XOR_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1202 gnd S0 addersubtractor_0/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1203 vdd S0 addersubtractor_0/XOR_0/NAND_2/in1 addersubtractor_0/XOR_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1204 addersubtractor_0/XOR_0/NAND_3/in1 enableblock_0/A_out2 addersubtractor_0/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1205 addersubtractor_0/XOR_0/NAND_3/in1 enableblock_0/A_out2 vdd addersubtractor_0/XOR_0/NAND_1/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1206 gnd addersubtractor_0/XOR_0/NAND_2/in1 addersubtractor_0/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1207 vdd addersubtractor_0/XOR_0/NAND_2/in1 addersubtractor_0/XOR_0/NAND_3/in1 addersubtractor_0/XOR_0/NAND_1/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1208 addersubtractor_0/XOR_0/NAND_3/in2 addersubtractor_0/XOR_0/NAND_2/in1 addersubtractor_0/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1209 addersubtractor_0/XOR_0/NAND_3/in2 addersubtractor_0/XOR_0/NAND_2/in1 vdd addersubtractor_0/XOR_0/NAND_2/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1210 gnd S0 addersubtractor_0/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1211 vdd S0 addersubtractor_0/XOR_0/NAND_3/in2 addersubtractor_0/XOR_0/NAND_2/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1212 addersubtractor_0/XOR_0/out addersubtractor_0/XOR_0/NAND_3/in1 addersubtractor_0/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1213 addersubtractor_0/XOR_0/out addersubtractor_0/XOR_0/NAND_3/in1 vdd addersubtractor_0/XOR_0/NAND_3/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1214 gnd addersubtractor_0/XOR_0/NAND_3/in2 addersubtractor_0/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1215 vdd addersubtractor_0/XOR_0/NAND_3/in2 addersubtractor_0/XOR_0/out addersubtractor_0/XOR_0/NAND_3/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1216 addersubtractor_0/XOR_1/NAND_2/in1 enableblock_0/A_out0 addersubtractor_0/XOR_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1217 addersubtractor_0/XOR_1/NAND_2/in1 enableblock_0/A_out0 vdd addersubtractor_0/XOR_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1218 gnd S0 addersubtractor_0/XOR_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1219 vdd S0 addersubtractor_0/XOR_1/NAND_2/in1 addersubtractor_0/XOR_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1220 addersubtractor_0/XOR_1/NAND_3/in1 enableblock_0/A_out0 addersubtractor_0/XOR_1/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1221 addersubtractor_0/XOR_1/NAND_3/in1 enableblock_0/A_out0 vdd addersubtractor_0/XOR_1/NAND_1/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1222 gnd addersubtractor_0/XOR_1/NAND_2/in1 addersubtractor_0/XOR_1/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1223 vdd addersubtractor_0/XOR_1/NAND_2/in1 addersubtractor_0/XOR_1/NAND_3/in1 addersubtractor_0/XOR_1/NAND_1/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1224 addersubtractor_0/XOR_1/NAND_3/in2 addersubtractor_0/XOR_1/NAND_2/in1 addersubtractor_0/XOR_1/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1225 addersubtractor_0/XOR_1/NAND_3/in2 addersubtractor_0/XOR_1/NAND_2/in1 vdd addersubtractor_0/XOR_1/NAND_2/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1226 gnd S0 addersubtractor_0/XOR_1/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1227 vdd S0 addersubtractor_0/XOR_1/NAND_3/in2 addersubtractor_0/XOR_1/NAND_2/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1228 addersubtractor_0/XOR_1/out addersubtractor_0/XOR_1/NAND_3/in1 addersubtractor_0/XOR_1/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1229 addersubtractor_0/XOR_1/out addersubtractor_0/XOR_1/NAND_3/in1 vdd addersubtractor_0/XOR_1/NAND_3/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1230 gnd addersubtractor_0/XOR_1/NAND_3/in2 addersubtractor_0/XOR_1/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1231 vdd addersubtractor_0/XOR_1/NAND_3/in2 addersubtractor_0/XOR_1/out addersubtractor_0/XOR_1/NAND_3/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1232 addersubtractor_0/XOR_2/NAND_2/in1 enableblock_0/B_out2 addersubtractor_0/XOR_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1233 addersubtractor_0/XOR_2/NAND_2/in1 enableblock_0/B_out2 vdd addersubtractor_0/XOR_2/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1234 gnd S0 addersubtractor_0/XOR_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1235 vdd S0 addersubtractor_0/XOR_2/NAND_2/in1 addersubtractor_0/XOR_2/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1236 addersubtractor_0/XOR_2/NAND_3/in1 enableblock_0/B_out2 addersubtractor_0/XOR_2/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1237 addersubtractor_0/XOR_2/NAND_3/in1 enableblock_0/B_out2 vdd addersubtractor_0/XOR_2/NAND_1/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1238 gnd addersubtractor_0/XOR_2/NAND_2/in1 addersubtractor_0/XOR_2/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1239 vdd addersubtractor_0/XOR_2/NAND_2/in1 addersubtractor_0/XOR_2/NAND_3/in1 addersubtractor_0/XOR_2/NAND_1/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1240 addersubtractor_0/XOR_2/NAND_3/in2 addersubtractor_0/XOR_2/NAND_2/in1 addersubtractor_0/XOR_2/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1241 addersubtractor_0/XOR_2/NAND_3/in2 addersubtractor_0/XOR_2/NAND_2/in1 vdd addersubtractor_0/XOR_2/NAND_2/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1242 gnd S0 addersubtractor_0/XOR_2/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1243 vdd S0 addersubtractor_0/XOR_2/NAND_3/in2 addersubtractor_0/XOR_2/NAND_2/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1244 addersubtractor_0/XOR_2/out addersubtractor_0/XOR_2/NAND_3/in1 addersubtractor_0/XOR_2/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1245 addersubtractor_0/XOR_2/out addersubtractor_0/XOR_2/NAND_3/in1 vdd addersubtractor_0/XOR_2/NAND_3/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1246 gnd addersubtractor_0/XOR_2/NAND_3/in2 addersubtractor_0/XOR_2/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1247 vdd addersubtractor_0/XOR_2/NAND_3/in2 addersubtractor_0/XOR_2/out addersubtractor_0/XOR_2/NAND_3/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1248 addersubtractor_0/XOR_3/NAND_2/in1 enableblock_0/B_out0 addersubtractor_0/XOR_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1249 addersubtractor_0/XOR_3/NAND_2/in1 enableblock_0/B_out0 vdd addersubtractor_0/XOR_3/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1250 gnd S0 addersubtractor_0/XOR_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1251 vdd S0 addersubtractor_0/XOR_3/NAND_2/in1 addersubtractor_0/XOR_3/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1252 addersubtractor_0/XOR_3/NAND_3/in1 enableblock_0/B_out0 addersubtractor_0/XOR_3/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1253 addersubtractor_0/XOR_3/NAND_3/in1 enableblock_0/B_out0 vdd addersubtractor_0/XOR_3/NAND_1/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1254 gnd addersubtractor_0/XOR_3/NAND_2/in1 addersubtractor_0/XOR_3/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1255 vdd addersubtractor_0/XOR_3/NAND_2/in1 addersubtractor_0/XOR_3/NAND_3/in1 addersubtractor_0/XOR_3/NAND_1/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1256 addersubtractor_0/XOR_3/NAND_3/in2 addersubtractor_0/XOR_3/NAND_2/in1 addersubtractor_0/XOR_3/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1257 addersubtractor_0/XOR_3/NAND_3/in2 addersubtractor_0/XOR_3/NAND_2/in1 vdd addersubtractor_0/XOR_3/NAND_2/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1258 gnd S0 addersubtractor_0/XOR_3/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1259 vdd S0 addersubtractor_0/XOR_3/NAND_3/in2 addersubtractor_0/XOR_3/NAND_2/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1260 addersubtractor_0/XOR_3/out addersubtractor_0/XOR_3/NAND_3/in1 addersubtractor_0/XOR_3/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1261 addersubtractor_0/XOR_3/out addersubtractor_0/XOR_3/NAND_3/in1 vdd addersubtractor_0/XOR_3/NAND_3/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1262 gnd addersubtractor_0/XOR_3/NAND_3/in2 addersubtractor_0/XOR_3/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1263 vdd addersubtractor_0/XOR_3/NAND_3/in2 addersubtractor_0/XOR_3/out addersubtractor_0/XOR_3/NAND_3/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1264 AND_0/not_0/in AND_0/in1 AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1265 AND_0/not_0/in AND_0/in1 vdd AND_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1266 gnd OR_0/out AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1267 vdd OR_0/out AND_0/not_0/in AND_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1268 XOR_0/in1 AND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1269 XOR_0/in1 AND_0/not_0/in vdd AND_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1270 AND_2/not_0/in AND_2/in1 AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1271 AND_2/not_0/in AND_2/in1 vdd AND_2/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1272 gnd AND_2/in2 AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1273 vdd AND_2/in2 AND_2/not_0/in AND_2/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1274 equal AND_2/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1275 equal AND_2/not_0/in vdd AND_2/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1276 enableblock_1/enable1_0/AND_0/not_0/in A3 enableblock_1/enable1_0/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1277 enableblock_1/enable1_0/AND_0/not_0/in A3 vdd enableblock_1/enable1_0/AND_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1278 gnd AND_2/in2 enableblock_1/enable1_0/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1279 vdd AND_2/in2 enableblock_1/enable1_0/AND_0/not_0/in enableblock_1/enable1_0/AND_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1280 comparator_0/A3 enableblock_1/enable1_0/AND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1281 comparator_0/A3 enableblock_1/enable1_0/AND_0/not_0/in vdd enableblock_1/enable1_0/AND_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1282 enableblock_1/enable1_0/AND_1/not_0/in AND_2/in2 enableblock_1/enable1_0/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1283 enableblock_1/enable1_0/AND_1/not_0/in AND_2/in2 vdd enableblock_1/enable1_0/AND_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1284 gnd B3 enableblock_1/enable1_0/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1285 vdd B3 enableblock_1/enable1_0/AND_1/not_0/in enableblock_1/enable1_0/AND_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1286 comparator_0/B3 enableblock_1/enable1_0/AND_1/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1287 comparator_0/B3 enableblock_1/enable1_0/AND_1/not_0/in vdd enableblock_1/enable1_0/AND_1/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1288 enableblock_1/enable1_0/AND_2/not_0/in A2 enableblock_1/enable1_0/AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1289 enableblock_1/enable1_0/AND_2/not_0/in A2 vdd enableblock_1/enable1_0/AND_2/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1290 gnd AND_2/in2 enableblock_1/enable1_0/AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1291 vdd AND_2/in2 enableblock_1/enable1_0/AND_2/not_0/in enableblock_1/enable1_0/AND_2/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1292 comparator_0/A2 enableblock_1/enable1_0/AND_2/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1293 comparator_0/A2 enableblock_1/enable1_0/AND_2/not_0/in vdd enableblock_1/enable1_0/AND_2/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1294 enableblock_1/enable1_0/AND_3/not_0/in AND_2/in2 enableblock_1/enable1_0/AND_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1295 enableblock_1/enable1_0/AND_3/not_0/in AND_2/in2 vdd enableblock_1/enable1_0/AND_3/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1296 gnd B2 enableblock_1/enable1_0/AND_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1297 vdd B2 enableblock_1/enable1_0/AND_3/not_0/in enableblock_1/enable1_0/AND_3/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1298 comparator_0/B2 enableblock_1/enable1_0/AND_3/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1299 comparator_0/B2 enableblock_1/enable1_0/AND_3/not_0/in vdd enableblock_1/enable1_0/AND_3/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1300 enableblock_1/enable1_1/AND_0/not_0/in A1 enableblock_1/enable1_1/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1301 enableblock_1/enable1_1/AND_0/not_0/in A1 vdd enableblock_1/enable1_1/AND_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1302 gnd AND_2/in2 enableblock_1/enable1_1/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1303 vdd AND_2/in2 enableblock_1/enable1_1/AND_0/not_0/in enableblock_1/enable1_1/AND_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1304 comparator_0/A1 enableblock_1/enable1_1/AND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1305 comparator_0/A1 enableblock_1/enable1_1/AND_0/not_0/in vdd enableblock_1/enable1_1/AND_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1306 enableblock_1/enable1_1/AND_1/not_0/in AND_2/in2 enableblock_1/enable1_1/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1307 enableblock_1/enable1_1/AND_1/not_0/in AND_2/in2 vdd enableblock_1/enable1_1/AND_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1308 gnd B1 enableblock_1/enable1_1/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1309 vdd B1 enableblock_1/enable1_1/AND_1/not_0/in enableblock_1/enable1_1/AND_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1310 comparator_0/B1 enableblock_1/enable1_1/AND_1/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1311 comparator_0/B1 enableblock_1/enable1_1/AND_1/not_0/in vdd enableblock_1/enable1_1/AND_1/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1312 enableblock_1/enable1_1/AND_2/not_0/in A0 enableblock_1/enable1_1/AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1313 enableblock_1/enable1_1/AND_2/not_0/in A0 vdd enableblock_1/enable1_1/AND_2/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1314 gnd AND_2/in2 enableblock_1/enable1_1/AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1315 vdd AND_2/in2 enableblock_1/enable1_1/AND_2/not_0/in enableblock_1/enable1_1/AND_2/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1316 comparator_0/A0 enableblock_1/enable1_1/AND_2/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1317 comparator_0/A0 enableblock_1/enable1_1/AND_2/not_0/in vdd enableblock_1/enable1_1/AND_2/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1318 enableblock_1/enable1_1/AND_3/not_0/in AND_2/in2 enableblock_1/enable1_1/AND_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1319 enableblock_1/enable1_1/AND_3/not_0/in AND_2/in2 vdd enableblock_1/enable1_1/AND_3/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1320 gnd B0 enableblock_1/enable1_1/AND_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1321 vdd B0 enableblock_1/enable1_1/AND_3/not_0/in enableblock_1/enable1_1/AND_3/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1322 comparator_0/B0 enableblock_1/enable1_1/AND_3/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1323 comparator_0/B0 enableblock_1/enable1_1/AND_3/not_0/in vdd enableblock_1/enable1_1/AND_3/not_0/w_0_0# CMOSP w=4 l=2
+  ad=45 pd=38 as=0 ps=0
M1324 enableblock_0/enable1_0/AND_0/not_0/in A0 enableblock_0/enable1_0/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1325 enableblock_0/enable1_0/AND_0/not_0/in A0 vdd enableblock_0/enable1_0/AND_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1326 gnd OR_0/out enableblock_0/enable1_0/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1327 vdd OR_0/out enableblock_0/enable1_0/AND_0/not_0/in enableblock_0/enable1_0/AND_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1328 enableblock_0/A_out3 enableblock_0/enable1_0/AND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1329 enableblock_0/A_out3 enableblock_0/enable1_0/AND_0/not_0/in vdd enableblock_0/enable1_0/AND_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1330 enableblock_0/enable1_0/AND_1/not_0/in OR_0/out enableblock_0/enable1_0/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1331 enableblock_0/enable1_0/AND_1/not_0/in OR_0/out vdd enableblock_0/enable1_0/AND_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1332 gnd B0 enableblock_0/enable1_0/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1333 vdd B0 enableblock_0/enable1_0/AND_1/not_0/in enableblock_0/enable1_0/AND_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1334 enableblock_0/A_out2 enableblock_0/enable1_0/AND_1/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1335 enableblock_0/A_out2 enableblock_0/enable1_0/AND_1/not_0/in vdd enableblock_0/enable1_0/AND_1/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1336 enableblock_0/enable1_0/AND_2/not_0/in A1 enableblock_0/enable1_0/AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1337 enableblock_0/enable1_0/AND_2/not_0/in A1 vdd enableblock_0/enable1_0/AND_2/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1338 gnd OR_0/out enableblock_0/enable1_0/AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1339 vdd OR_0/out enableblock_0/enable1_0/AND_2/not_0/in enableblock_0/enable1_0/AND_2/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1340 enableblock_0/A_out1 enableblock_0/enable1_0/AND_2/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1341 enableblock_0/A_out1 enableblock_0/enable1_0/AND_2/not_0/in vdd enableblock_0/enable1_0/AND_2/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1342 enableblock_0/enable1_0/AND_3/not_0/in OR_0/out enableblock_0/enable1_0/AND_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1343 enableblock_0/enable1_0/AND_3/not_0/in OR_0/out vdd enableblock_0/enable1_0/AND_3/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1344 gnd B1 enableblock_0/enable1_0/AND_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1345 vdd B1 enableblock_0/enable1_0/AND_3/not_0/in enableblock_0/enable1_0/AND_3/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1346 enableblock_0/A_out0 enableblock_0/enable1_0/AND_3/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1347 enableblock_0/A_out0 enableblock_0/enable1_0/AND_3/not_0/in vdd enableblock_0/enable1_0/AND_3/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1348 enableblock_0/enable1_1/AND_0/not_0/in A2 enableblock_0/enable1_1/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1349 enableblock_0/enable1_1/AND_0/not_0/in A2 vdd enableblock_0/enable1_1/AND_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1350 gnd OR_0/out enableblock_0/enable1_1/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1351 vdd OR_0/out enableblock_0/enable1_1/AND_0/not_0/in enableblock_0/enable1_1/AND_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1352 enableblock_0/B_out3 enableblock_0/enable1_1/AND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1353 enableblock_0/B_out3 enableblock_0/enable1_1/AND_0/not_0/in vdd enableblock_0/enable1_1/AND_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1354 enableblock_0/enable1_1/AND_1/not_0/in OR_0/out enableblock_0/enable1_1/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1355 enableblock_0/enable1_1/AND_1/not_0/in OR_0/out vdd enableblock_0/enable1_1/AND_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1356 gnd B2 enableblock_0/enable1_1/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1357 vdd B2 enableblock_0/enable1_1/AND_1/not_0/in enableblock_0/enable1_1/AND_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1358 enableblock_0/B_out2 enableblock_0/enable1_1/AND_1/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1359 enableblock_0/B_out2 enableblock_0/enable1_1/AND_1/not_0/in vdd enableblock_0/enable1_1/AND_1/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1360 enableblock_0/enable1_1/AND_2/not_0/in A3 enableblock_0/enable1_1/AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1361 enableblock_0/enable1_1/AND_2/not_0/in A3 vdd enableblock_0/enable1_1/AND_2/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1362 gnd OR_0/out enableblock_0/enable1_1/AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1363 vdd OR_0/out enableblock_0/enable1_1/AND_2/not_0/in enableblock_0/enable1_1/AND_2/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1364 enableblock_0/B_out1 enableblock_0/enable1_1/AND_2/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1365 enableblock_0/B_out1 enableblock_0/enable1_1/AND_2/not_0/in vdd enableblock_0/enable1_1/AND_2/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1366 enableblock_0/enable1_1/AND_3/not_0/in OR_0/out enableblock_0/enable1_1/AND_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1367 enableblock_0/enable1_1/AND_3/not_0/in OR_0/out vdd enableblock_0/enable1_1/AND_3/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1368 gnd B3 enableblock_0/enable1_1/AND_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1369 vdd B3 enableblock_0/enable1_1/AND_3/not_0/in enableblock_0/enable1_1/AND_3/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1370 enableblock_0/B_out0 enableblock_0/enable1_1/AND_3/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1371 enableblock_0/B_out0 enableblock_0/enable1_1/AND_3/not_0/in vdd enableblock_0/enable1_1/AND_3/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1372 enableblock_2/enable1_0/AND_0/not_0/in A3 enableblock_2/enable1_0/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1373 enableblock_2/enable1_0/AND_0/not_0/in A3 vdd enableblock_2/enable1_0/AND_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1374 gnd enableblock_2/En enableblock_2/enable1_0/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1375 vdd enableblock_2/En enableblock_2/enable1_0/AND_0/not_0/in enableblock_2/enable1_0/AND_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1376 andblock_0/A3 enableblock_2/enable1_0/AND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1377 andblock_0/A3 enableblock_2/enable1_0/AND_0/not_0/in vdd enableblock_2/enable1_0/AND_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1378 enableblock_2/enable1_0/AND_1/not_0/in enableblock_2/En enableblock_2/enable1_0/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1379 enableblock_2/enable1_0/AND_1/not_0/in enableblock_2/En vdd enableblock_2/enable1_0/AND_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1380 gnd B3 enableblock_2/enable1_0/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1381 vdd B3 enableblock_2/enable1_0/AND_1/not_0/in enableblock_2/enable1_0/AND_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1382 andblock_0/B3 enableblock_2/enable1_0/AND_1/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1383 andblock_0/B3 enableblock_2/enable1_0/AND_1/not_0/in vdd enableblock_2/enable1_0/AND_1/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1384 enableblock_2/enable1_0/AND_2/not_0/in A2 enableblock_2/enable1_0/AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1385 enableblock_2/enable1_0/AND_2/not_0/in A2 vdd enableblock_2/enable1_0/AND_2/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1386 gnd enableblock_2/En enableblock_2/enable1_0/AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1387 vdd enableblock_2/En enableblock_2/enable1_0/AND_2/not_0/in enableblock_2/enable1_0/AND_2/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1388 andblock_0/A2 enableblock_2/enable1_0/AND_2/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1389 andblock_0/A2 enableblock_2/enable1_0/AND_2/not_0/in vdd enableblock_2/enable1_0/AND_2/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1390 enableblock_2/enable1_0/AND_3/not_0/in enableblock_2/En enableblock_2/enable1_0/AND_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1391 enableblock_2/enable1_0/AND_3/not_0/in enableblock_2/En vdd enableblock_2/enable1_0/AND_3/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1392 gnd B2 enableblock_2/enable1_0/AND_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1393 vdd B2 enableblock_2/enable1_0/AND_3/not_0/in enableblock_2/enable1_0/AND_3/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1394 andblock_0/B2 enableblock_2/enable1_0/AND_3/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1395 andblock_0/B2 enableblock_2/enable1_0/AND_3/not_0/in vdd enableblock_2/enable1_0/AND_3/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1396 enableblock_2/enable1_1/AND_0/not_0/in A1 enableblock_2/enable1_1/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1397 enableblock_2/enable1_1/AND_0/not_0/in A1 vdd enableblock_2/enable1_1/AND_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1398 gnd enableblock_2/En enableblock_2/enable1_1/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1399 vdd enableblock_2/En enableblock_2/enable1_1/AND_0/not_0/in enableblock_2/enable1_1/AND_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1400 andblock_0/A1 enableblock_2/enable1_1/AND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1401 andblock_0/A1 enableblock_2/enable1_1/AND_0/not_0/in vdd enableblock_2/enable1_1/AND_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1402 enableblock_2/enable1_1/AND_1/not_0/in enableblock_2/En enableblock_2/enable1_1/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1403 enableblock_2/enable1_1/AND_1/not_0/in enableblock_2/En vdd enableblock_2/enable1_1/AND_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1404 gnd B1 enableblock_2/enable1_1/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1405 vdd B1 enableblock_2/enable1_1/AND_1/not_0/in enableblock_2/enable1_1/AND_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1406 andblock_0/B1 enableblock_2/enable1_1/AND_1/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1407 andblock_0/B1 enableblock_2/enable1_1/AND_1/not_0/in vdd enableblock_2/enable1_1/AND_1/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1408 enableblock_2/enable1_1/AND_2/not_0/in A0 enableblock_2/enable1_1/AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1409 enableblock_2/enable1_1/AND_2/not_0/in A0 vdd enableblock_2/enable1_1/AND_2/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1410 gnd enableblock_2/En enableblock_2/enable1_1/AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1411 vdd enableblock_2/En enableblock_2/enable1_1/AND_2/not_0/in enableblock_2/enable1_1/AND_2/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1412 andblock_0/A0 enableblock_2/enable1_1/AND_2/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1413 andblock_0/A0 enableblock_2/enable1_1/AND_2/not_0/in vdd enableblock_2/enable1_1/AND_2/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1414 enableblock_2/enable1_1/AND_3/not_0/in enableblock_2/En enableblock_2/enable1_1/AND_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1415 enableblock_2/enable1_1/AND_3/not_0/in enableblock_2/En vdd enableblock_2/enable1_1/AND_3/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1416 gnd B0 enableblock_2/enable1_1/AND_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1417 vdd B0 enableblock_2/enable1_1/AND_3/not_0/in enableblock_2/enable1_1/AND_3/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1418 andblock_0/B0 enableblock_2/enable1_1/AND_3/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1419 andblock_0/B0 enableblock_2/enable1_1/AND_3/not_0/in vdd enableblock_2/enable1_1/AND_3/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1420 twotofourdecoder_0/AND_0/not_0/in S0 twotofourdecoder_0/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1421 twotofourdecoder_0/AND_0/not_0/in S0 vdd twotofourdecoder_0/AND_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1422 gnd S1 twotofourdecoder_0/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1423 vdd S1 twotofourdecoder_0/AND_0/not_0/in twotofourdecoder_0/AND_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1424 enableblock_2/En twotofourdecoder_0/AND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1425 enableblock_2/En twotofourdecoder_0/AND_0/not_0/in vdd twotofourdecoder_0/AND_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1426 twotofourdecoder_0/AND_1/not_0/in S1 twotofourdecoder_0/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1427 twotofourdecoder_0/AND_1/not_0/in S1 vdd twotofourdecoder_0/AND_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1428 gnd twotofourdecoder_0/not_0/out twotofourdecoder_0/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1429 vdd twotofourdecoder_0/not_0/out twotofourdecoder_0/AND_1/not_0/in twotofourdecoder_0/AND_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1430 AND_2/in2 twotofourdecoder_0/AND_1/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1431 AND_2/in2 twotofourdecoder_0/AND_1/not_0/in vdd twotofourdecoder_0/AND_1/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1432 twotofourdecoder_0/AND_2/not_0/in twotofourdecoder_0/not_0/out twotofourdecoder_0/AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1433 twotofourdecoder_0/AND_2/not_0/in twotofourdecoder_0/not_0/out vdd twotofourdecoder_0/AND_2/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1434 gnd twotofourdecoder_0/not_1/out twotofourdecoder_0/AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1435 vdd twotofourdecoder_0/not_1/out twotofourdecoder_0/AND_2/not_0/in twotofourdecoder_0/AND_2/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1436 OR_0/in2 twotofourdecoder_0/AND_2/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1437 OR_0/in2 twotofourdecoder_0/AND_2/not_0/in vdd twotofourdecoder_0/AND_2/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1438 twotofourdecoder_0/AND_3/not_0/in twotofourdecoder_0/not_1/out twotofourdecoder_0/AND_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1439 twotofourdecoder_0/AND_3/not_0/in twotofourdecoder_0/not_1/out vdd twotofourdecoder_0/AND_3/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1440 gnd S0 twotofourdecoder_0/AND_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1441 vdd S0 twotofourdecoder_0/AND_3/not_0/in twotofourdecoder_0/AND_3/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1442 OR_0/in1 twotofourdecoder_0/AND_3/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1443 OR_0/in1 twotofourdecoder_0/AND_3/not_0/in vdd twotofourdecoder_0/AND_3/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1444 twotofourdecoder_0/not_0/out S0 gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1445 twotofourdecoder_0/not_0/out S0 vdd twotofourdecoder_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1446 twotofourdecoder_0/not_1/out S1 gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1447 twotofourdecoder_0/not_1/out S1 vdd twotofourdecoder_0/not_1/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1448 comparator_0/fourinputOR_0/not_0/in comparator_0/fourinputOR_0/in4 gnd Gnd CMOSN w=4 l=2
+  ad=80 pd=72 as=0 ps=0
M1449 comparator_0/fourinputOR_0/not_0/in comparator_0/AND_0/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1450 comparator_0/fourinputOR_0/fourinputNOR_0/a_77_6# comparator_0/fourinputOR_0/in3 comparator_0/fourinputOR_0/fourinputNOR_0/a_45_6# comparator_0/fourinputOR_0/fourinputNOR_0/w_64_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=40 ps=36
M1451 comparator_0/fourinputOR_0/not_0/in comparator_0/fourinputOR_0/in3 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1452 comparator_0/fourinputOR_0/fourinputNOR_0/a_13_6# comparator_0/AND_0/out vdd comparator_0/fourinputOR_0/fourinputNOR_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1453 comparator_0/fourinputOR_0/not_0/in comparator_0/fourinputOR_0/in4 comparator_0/fourinputOR_0/fourinputNOR_0/a_77_6# comparator_0/fourinputOR_0/fourinputNOR_0/w_97_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1454 gnd comparator_0/fourinputOR_0/in2 comparator_0/fourinputOR_0/not_0/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1455 comparator_0/fourinputOR_0/fourinputNOR_0/a_45_6# comparator_0/fourinputOR_0/in2 comparator_0/fourinputOR_0/fourinputNOR_0/a_13_6# comparator_0/fourinputOR_0/fourinputNOR_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1456 greater comparator_0/fourinputOR_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1457 greater comparator_0/fourinputOR_0/not_0/in vdd comparator_0/fourinputOR_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1458 comparator_0/AND_0/not_0/in comparator_0/not_0/out comparator_0/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1459 comparator_0/AND_0/not_0/in comparator_0/not_0/out vdd comparator_0/AND_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1460 gnd comparator_0/A3 comparator_0/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1461 vdd comparator_0/A3 comparator_0/AND_0/not_0/in comparator_0/AND_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1462 comparator_0/AND_0/out comparator_0/AND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1463 comparator_0/AND_0/out comparator_0/AND_0/not_0/in vdd comparator_0/AND_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1464 comparator_0/not_0/out comparator_0/B3 gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1465 comparator_0/not_0/out comparator_0/B3 vdd comparator_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1466 comparator_0/not_1/out comparator_0/B2 gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1467 comparator_0/not_1/out comparator_0/B2 vdd comparator_0/not_1/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1468 comparator_0/not_2/out comparator_0/B1 gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1469 comparator_0/not_2/out comparator_0/B1 vdd comparator_0/not_2/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1470 comparator_0/not_3/out comparator_0/B0 gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1471 comparator_0/not_3/out comparator_0/B0 vdd comparator_0/not_3/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1472 comparator_0/fourinputOR_0/in3 comparator_0/fourinputAND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1473 comparator_0/fourinputOR_0/in3 comparator_0/fourinputAND_0/not_0/in vdd comparator_0/fourinputAND_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1474 comparator_0/fourinputAND_0/not_0/in comparator_0/not_2/out comparator_0/fourinputAND_0/fourinputNAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1475 gnd comparator_0/XNOR_0/out comparator_0/fourinputAND_0/fourinputNAND_0/a_76_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1476 comparator_0/fourinputAND_0/not_0/in comparator_0/XNOR_1/out vdd comparator_0/fourinputAND_0/fourinputNAND_0/w_63_0# CMOSP w=4 l=2
+  ad=80 pd=72 as=0 ps=0
M1477 comparator_0/fourinputAND_0/not_0/in comparator_0/not_2/out vdd comparator_0/fourinputAND_0/fourinputNAND_0/w_0_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1478 comparator_0/fourinputAND_0/fourinputNAND_0/a_76_n14# comparator_0/XNOR_1/out comparator_0/fourinputAND_0/fourinputNAND_0/a_45_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1479 comparator_0/fourinputAND_0/fourinputNAND_0/a_45_n14# comparator_0/A1 comparator_0/fourinputAND_0/fourinputNAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1480 vdd comparator_0/A1 comparator_0/fourinputAND_0/not_0/in comparator_0/fourinputAND_0/fourinputNAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1481 vdd comparator_0/XNOR_0/out comparator_0/fourinputAND_0/not_0/in comparator_0/fourinputAND_0/fourinputNAND_0/w_100_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1482 AND_2/in1 comparator_0/fourinputAND_1/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1483 AND_2/in1 comparator_0/fourinputAND_1/not_0/in vdd comparator_0/fourinputAND_1/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1484 comparator_0/fourinputAND_1/not_0/in comparator_0/XNOR_3/out comparator_0/fourinputAND_1/fourinputNAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1485 gnd comparator_0/XNOR_2/out comparator_0/fourinputAND_1/fourinputNAND_0/a_76_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1486 comparator_0/fourinputAND_1/not_0/in comparator_0/XNOR_1/out vdd comparator_0/fourinputAND_1/fourinputNAND_0/w_63_0# CMOSP w=4 l=2
+  ad=80 pd=72 as=0 ps=0
M1487 comparator_0/fourinputAND_1/not_0/in comparator_0/XNOR_3/out vdd comparator_0/fourinputAND_1/fourinputNAND_0/w_0_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1488 comparator_0/fourinputAND_1/fourinputNAND_0/a_76_n14# comparator_0/XNOR_1/out comparator_0/fourinputAND_1/fourinputNAND_0/a_45_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1489 comparator_0/fourinputAND_1/fourinputNAND_0/a_45_n14# comparator_0/XNOR_0/out comparator_0/fourinputAND_1/fourinputNAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1490 vdd comparator_0/XNOR_0/out comparator_0/fourinputAND_1/not_0/in comparator_0/fourinputAND_1/fourinputNAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1491 vdd comparator_0/XNOR_2/out comparator_0/fourinputAND_1/not_0/in comparator_0/fourinputAND_1/fourinputNAND_0/w_100_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1492 comparator_0/threeinputAND_0/not_0/in comparator_0/not_1/out comparator_0/threeinputAND_0/threeinputNAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1493 comparator_0/threeinputAND_0/not_0/in comparator_0/XNOR_0/out vdd comparator_0/threeinputAND_0/threeinputNAND_0/w_63_0# CMOSP w=4 l=2
+  ad=60 pd=54 as=0 ps=0
M1494 comparator_0/threeinputAND_0/not_0/in comparator_0/not_1/out vdd comparator_0/threeinputAND_0/threeinputNAND_0/w_0_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1495 gnd comparator_0/XNOR_0/out comparator_0/threeinputAND_0/threeinputNAND_0/a_45_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1496 comparator_0/threeinputAND_0/threeinputNAND_0/a_45_n14# comparator_0/A2 comparator_0/threeinputAND_0/threeinputNAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1497 vdd comparator_0/A2 comparator_0/threeinputAND_0/not_0/in comparator_0/threeinputAND_0/threeinputNAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1498 comparator_0/fourinputOR_0/in2 comparator_0/threeinputAND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1499 comparator_0/fourinputOR_0/in2 comparator_0/threeinputAND_0/not_0/in vdd comparator_0/threeinputAND_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1500 comparator_0/fourinputOR_0/in4 comparator_0/fiveinputAND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1501 comparator_0/fourinputOR_0/in4 comparator_0/fiveinputAND_0/not_0/in vdd comparator_0/fiveinputAND_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1502 comparator_0/fiveinputAND_0/not_0/in comparator_0/not_3/out comparator_0/fiveinputAND_0/fiveinputNAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1503 comparator_0/fiveinputAND_0/fiveinputNAND_0/a_113_n14# comparator_0/XNOR_0/out comparator_0/fiveinputAND_0/fiveinputNAND_0/a_76_n14# Gnd CMOSN w=4 l=2
+  ad=40 pd=36 as=40 ps=36
M1504 comparator_0/fiveinputAND_0/not_0/in comparator_0/XNOR_2/out vdd comparator_0/fiveinputAND_0/fiveinputNAND_0/w_133_0# CMOSP w=4 l=2
+  ad=100 pd=90 as=0 ps=0
M1505 comparator_0/fiveinputAND_0/not_0/in comparator_0/XNOR_1/out vdd comparator_0/fiveinputAND_0/fiveinputNAND_0/w_63_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1506 comparator_0/fiveinputAND_0/not_0/in comparator_0/not_3/out vdd comparator_0/fiveinputAND_0/fiveinputNAND_0/w_0_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1507 gnd comparator_0/XNOR_2/out comparator_0/fiveinputAND_0/fiveinputNAND_0/a_113_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1508 comparator_0/fiveinputAND_0/fiveinputNAND_0/a_76_n14# comparator_0/XNOR_1/out comparator_0/fiveinputAND_0/fiveinputNAND_0/a_45_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1509 comparator_0/fiveinputAND_0/fiveinputNAND_0/a_45_n14# comparator_0/A0 comparator_0/fiveinputAND_0/fiveinputNAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1510 vdd comparator_0/A0 comparator_0/fiveinputAND_0/not_0/in comparator_0/fiveinputAND_0/fiveinputNAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1511 vdd comparator_0/XNOR_0/out comparator_0/fiveinputAND_0/not_0/in comparator_0/fiveinputAND_0/fiveinputNAND_0/w_100_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1512 comparator_0/XNOR_1/out comparator_0/XNOR_1/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1513 comparator_0/XNOR_1/out comparator_0/XNOR_1/not_0/in vdd comparator_0/XNOR_1/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1514 comparator_0/XNOR_1/XOR_0/NAND_2/in1 comparator_0/A2 comparator_0/XNOR_1/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1515 comparator_0/XNOR_1/XOR_0/NAND_2/in1 comparator_0/A2 vdd comparator_0/XNOR_1/XOR_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1516 gnd comparator_0/B2 comparator_0/XNOR_1/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1517 vdd comparator_0/B2 comparator_0/XNOR_1/XOR_0/NAND_2/in1 comparator_0/XNOR_1/XOR_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1518 comparator_0/XNOR_1/XOR_0/NAND_3/in1 comparator_0/A2 comparator_0/XNOR_1/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1519 comparator_0/XNOR_1/XOR_0/NAND_3/in1 comparator_0/A2 vdd comparator_0/XNOR_1/XOR_0/NAND_1/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1520 gnd comparator_0/XNOR_1/XOR_0/NAND_2/in1 comparator_0/XNOR_1/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1521 vdd comparator_0/XNOR_1/XOR_0/NAND_2/in1 comparator_0/XNOR_1/XOR_0/NAND_3/in1 comparator_0/XNOR_1/XOR_0/NAND_1/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1522 comparator_0/XNOR_1/XOR_0/NAND_3/in2 comparator_0/XNOR_1/XOR_0/NAND_2/in1 comparator_0/XNOR_1/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1523 comparator_0/XNOR_1/XOR_0/NAND_3/in2 comparator_0/XNOR_1/XOR_0/NAND_2/in1 vdd comparator_0/XNOR_1/XOR_0/NAND_2/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1524 gnd comparator_0/B2 comparator_0/XNOR_1/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1525 vdd comparator_0/B2 comparator_0/XNOR_1/XOR_0/NAND_3/in2 comparator_0/XNOR_1/XOR_0/NAND_2/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1526 comparator_0/XNOR_1/not_0/in comparator_0/XNOR_1/XOR_0/NAND_3/in1 comparator_0/XNOR_1/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1527 comparator_0/XNOR_1/not_0/in comparator_0/XNOR_1/XOR_0/NAND_3/in1 vdd comparator_0/XNOR_1/XOR_0/NAND_3/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1528 gnd comparator_0/XNOR_1/XOR_0/NAND_3/in2 comparator_0/XNOR_1/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1529 vdd comparator_0/XNOR_1/XOR_0/NAND_3/in2 comparator_0/XNOR_1/not_0/in comparator_0/XNOR_1/XOR_0/NAND_3/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1530 comparator_0/XNOR_0/out comparator_0/XNOR_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1531 comparator_0/XNOR_0/out comparator_0/XNOR_0/not_0/in vdd comparator_0/XNOR_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1532 comparator_0/XNOR_0/XOR_0/NAND_2/in1 comparator_0/A3 comparator_0/XNOR_0/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1533 comparator_0/XNOR_0/XOR_0/NAND_2/in1 comparator_0/A3 vdd comparator_0/XNOR_0/XOR_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1534 gnd comparator_0/B3 comparator_0/XNOR_0/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1535 vdd comparator_0/B3 comparator_0/XNOR_0/XOR_0/NAND_2/in1 comparator_0/XNOR_0/XOR_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1536 comparator_0/XNOR_0/XOR_0/NAND_3/in1 comparator_0/A3 comparator_0/XNOR_0/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1537 comparator_0/XNOR_0/XOR_0/NAND_3/in1 comparator_0/A3 vdd comparator_0/XNOR_0/XOR_0/NAND_1/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1538 gnd comparator_0/XNOR_0/XOR_0/NAND_2/in1 comparator_0/XNOR_0/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1539 vdd comparator_0/XNOR_0/XOR_0/NAND_2/in1 comparator_0/XNOR_0/XOR_0/NAND_3/in1 comparator_0/XNOR_0/XOR_0/NAND_1/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1540 comparator_0/XNOR_0/XOR_0/NAND_3/in2 comparator_0/XNOR_0/XOR_0/NAND_2/in1 comparator_0/XNOR_0/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1541 comparator_0/XNOR_0/XOR_0/NAND_3/in2 comparator_0/XNOR_0/XOR_0/NAND_2/in1 vdd comparator_0/XNOR_0/XOR_0/NAND_2/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1542 gnd comparator_0/B3 comparator_0/XNOR_0/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1543 vdd comparator_0/B3 comparator_0/XNOR_0/XOR_0/NAND_3/in2 comparator_0/XNOR_0/XOR_0/NAND_2/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1544 comparator_0/XNOR_0/not_0/in comparator_0/XNOR_0/XOR_0/NAND_3/in1 comparator_0/XNOR_0/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1545 comparator_0/XNOR_0/not_0/in comparator_0/XNOR_0/XOR_0/NAND_3/in1 vdd comparator_0/XNOR_0/XOR_0/NAND_3/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1546 gnd comparator_0/XNOR_0/XOR_0/NAND_3/in2 comparator_0/XNOR_0/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1547 vdd comparator_0/XNOR_0/XOR_0/NAND_3/in2 comparator_0/XNOR_0/not_0/in comparator_0/XNOR_0/XOR_0/NAND_3/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1548 comparator_0/XNOR_2/out comparator_0/XNOR_2/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1549 comparator_0/XNOR_2/out comparator_0/XNOR_2/not_0/in vdd comparator_0/XNOR_2/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1550 comparator_0/XNOR_2/XOR_0/NAND_2/in1 comparator_0/A1 comparator_0/XNOR_2/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1551 comparator_0/XNOR_2/XOR_0/NAND_2/in1 comparator_0/A1 vdd comparator_0/XNOR_2/XOR_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1552 gnd comparator_0/B1 comparator_0/XNOR_2/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1553 vdd comparator_0/B1 comparator_0/XNOR_2/XOR_0/NAND_2/in1 comparator_0/XNOR_2/XOR_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1554 comparator_0/XNOR_2/XOR_0/NAND_3/in1 comparator_0/A1 comparator_0/XNOR_2/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1555 comparator_0/XNOR_2/XOR_0/NAND_3/in1 comparator_0/A1 vdd comparator_0/XNOR_2/XOR_0/NAND_1/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1556 gnd comparator_0/XNOR_2/XOR_0/NAND_2/in1 comparator_0/XNOR_2/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1557 vdd comparator_0/XNOR_2/XOR_0/NAND_2/in1 comparator_0/XNOR_2/XOR_0/NAND_3/in1 comparator_0/XNOR_2/XOR_0/NAND_1/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1558 comparator_0/XNOR_2/XOR_0/NAND_3/in2 comparator_0/XNOR_2/XOR_0/NAND_2/in1 comparator_0/XNOR_2/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1559 comparator_0/XNOR_2/XOR_0/NAND_3/in2 comparator_0/XNOR_2/XOR_0/NAND_2/in1 vdd comparator_0/XNOR_2/XOR_0/NAND_2/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1560 gnd comparator_0/B1 comparator_0/XNOR_2/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1561 vdd comparator_0/B1 comparator_0/XNOR_2/XOR_0/NAND_3/in2 comparator_0/XNOR_2/XOR_0/NAND_2/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1562 comparator_0/XNOR_2/not_0/in comparator_0/XNOR_2/XOR_0/NAND_3/in1 comparator_0/XNOR_2/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1563 comparator_0/XNOR_2/not_0/in comparator_0/XNOR_2/XOR_0/NAND_3/in1 vdd comparator_0/XNOR_2/XOR_0/NAND_3/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1564 gnd comparator_0/XNOR_2/XOR_0/NAND_3/in2 comparator_0/XNOR_2/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1565 vdd comparator_0/XNOR_2/XOR_0/NAND_3/in2 comparator_0/XNOR_2/not_0/in comparator_0/XNOR_2/XOR_0/NAND_3/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1566 comparator_0/XNOR_3/out comparator_0/XNOR_3/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1567 comparator_0/XNOR_3/out comparator_0/XNOR_3/not_0/in vdd comparator_0/XNOR_3/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1568 comparator_0/XNOR_3/XOR_0/NAND_2/in1 comparator_0/A0 comparator_0/XNOR_3/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1569 comparator_0/XNOR_3/XOR_0/NAND_2/in1 comparator_0/A0 vdd comparator_0/XNOR_3/XOR_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1570 gnd comparator_0/B0 comparator_0/XNOR_3/XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1571 vdd comparator_0/B0 comparator_0/XNOR_3/XOR_0/NAND_2/in1 comparator_0/XNOR_3/XOR_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1572 comparator_0/XNOR_3/XOR_0/NAND_3/in1 comparator_0/A0 comparator_0/XNOR_3/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1573 comparator_0/XNOR_3/XOR_0/NAND_3/in1 comparator_0/A0 vdd comparator_0/XNOR_3/XOR_0/NAND_1/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1574 gnd comparator_0/XNOR_3/XOR_0/NAND_2/in1 comparator_0/XNOR_3/XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1575 vdd comparator_0/XNOR_3/XOR_0/NAND_2/in1 comparator_0/XNOR_3/XOR_0/NAND_3/in1 comparator_0/XNOR_3/XOR_0/NAND_1/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1576 comparator_0/XNOR_3/XOR_0/NAND_3/in2 comparator_0/XNOR_3/XOR_0/NAND_2/in1 comparator_0/XNOR_3/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1577 comparator_0/XNOR_3/XOR_0/NAND_3/in2 comparator_0/XNOR_3/XOR_0/NAND_2/in1 vdd comparator_0/XNOR_3/XOR_0/NAND_2/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1578 gnd comparator_0/B0 comparator_0/XNOR_3/XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1579 vdd comparator_0/B0 comparator_0/XNOR_3/XOR_0/NAND_3/in2 comparator_0/XNOR_3/XOR_0/NAND_2/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1580 comparator_0/XNOR_3/not_0/in comparator_0/XNOR_3/XOR_0/NAND_3/in1 comparator_0/XNOR_3/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1581 comparator_0/XNOR_3/not_0/in comparator_0/XNOR_3/XOR_0/NAND_3/in1 vdd comparator_0/XNOR_3/XOR_0/NAND_3/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1582 gnd comparator_0/XNOR_3/XOR_0/NAND_3/in2 comparator_0/XNOR_3/XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1583 vdd comparator_0/XNOR_3/XOR_0/NAND_3/in2 comparator_0/XNOR_3/not_0/in comparator_0/XNOR_3/XOR_0/NAND_3/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1584 lesser greater gnd Gnd CMOSN w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1585 comparator_0/NOR_0/a_13_6# greater vdd comparator_0/NOR_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1586 gnd AND_2/in1 lesser Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1587 lesser AND_2/in1 comparator_0/NOR_0/a_13_6# comparator_0/NOR_0/w_32_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1588 andblock_0/AND_0/not_0/in andblock_0/A3 andblock_0/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1589 andblock_0/AND_0/not_0/in andblock_0/A3 vdd andblock_0/AND_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1590 gnd andblock_0/B3 andblock_0/AND_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1591 vdd andblock_0/B3 andblock_0/AND_0/not_0/in andblock_0/AND_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1592 and3 andblock_0/AND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1593 and3 andblock_0/AND_0/not_0/in vdd andblock_0/AND_0/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1594 andblock_0/AND_1/not_0/in andblock_0/A2 andblock_0/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1595 andblock_0/AND_1/not_0/in andblock_0/A2 vdd andblock_0/AND_1/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1596 gnd andblock_0/B2 andblock_0/AND_1/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1597 vdd andblock_0/B2 andblock_0/AND_1/not_0/in andblock_0/AND_1/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1598 and2 andblock_0/AND_1/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1599 and2 andblock_0/AND_1/not_0/in vdd andblock_0/AND_1/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1600 andblock_0/AND_2/not_0/in andblock_0/A1 andblock_0/AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1601 andblock_0/AND_2/not_0/in andblock_0/A1 vdd andblock_0/AND_2/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1602 gnd andblock_0/B1 andblock_0/AND_2/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1603 vdd andblock_0/B1 andblock_0/AND_2/not_0/in andblock_0/AND_2/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1604 and1 andblock_0/AND_2/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1605 and1 andblock_0/AND_2/not_0/in vdd andblock_0/AND_2/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1606 andblock_0/AND_3/not_0/in andblock_0/A0 andblock_0/AND_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1607 andblock_0/AND_3/not_0/in andblock_0/A0 vdd andblock_0/AND_3/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1608 gnd andblock_0/B0 andblock_0/AND_3/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1609 vdd andblock_0/B0 andblock_0/AND_3/not_0/in andblock_0/AND_3/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1610 and0 andblock_0/AND_3/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1611 and0 andblock_0/AND_3/not_0/in vdd andblock_0/AND_3/not_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1612 XOR_0/NAND_2/in1 XOR_0/in1 XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1613 XOR_0/NAND_2/in1 XOR_0/in1 vdd XOR_0/NAND_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1614 gnd OR_0/in1 XOR_0/NAND_0/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1615 vdd OR_0/in1 XOR_0/NAND_2/in1 XOR_0/NAND_0/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1616 XOR_0/NAND_3/in1 XOR_0/in1 XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1617 XOR_0/NAND_3/in1 XOR_0/in1 vdd XOR_0/NAND_1/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1618 gnd XOR_0/NAND_2/in1 XOR_0/NAND_1/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1619 vdd XOR_0/NAND_2/in1 XOR_0/NAND_3/in1 XOR_0/NAND_1/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1620 XOR_0/NAND_3/in2 XOR_0/NAND_2/in1 XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1621 XOR_0/NAND_3/in2 XOR_0/NAND_2/in1 vdd XOR_0/NAND_2/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1622 gnd OR_0/in1 XOR_0/NAND_2/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1623 vdd OR_0/in1 XOR_0/NAND_3/in2 XOR_0/NAND_2/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1624 Carry XOR_0/NAND_3/in1 XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1625 Carry XOR_0/NAND_3/in1 vdd XOR_0/NAND_3/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1626 gnd XOR_0/NAND_3/in2 XOR_0/NAND_3/a_6_n14# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1627 vdd XOR_0/NAND_3/in2 Carry XOR_0/NAND_3/w_32_0# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1628 OR_0/out OR_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1629 OR_0/out OR_0/NOT_0/in vdd OR_0/NOT_0/w_0_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1630 OR_0/NOT_0/in OR_0/in1 gnd Gnd CMOSN w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1631 OR_0/NOR_0/a_13_6# OR_0/in1 vdd OR_0/NOR_0/w_0_0# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1632 gnd OR_0/in2 OR_0/NOT_0/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1633 OR_0/NOT_0/in OR_0/in2 OR_0/NOR_0/a_13_6# OR_0/NOR_0/w_32_0# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
C0 AND_2/NAND_0/a_6_n14# AND_2/in1 0.08fF
C1 vdd comparator_0/XNOR_1/out 0.36fF
C2 AND_2/in2 enableblock_1/enable1_1/AND_0/NAND_0/w_32_0# 0.06fF
C3 enableblock_0/enable1_1/AND_1/NAND_0/w_32_0# B2 0.06fF
C4 gnd AND_2/in2 3.60fF
C5 addersubtractor_0/fulladder_2/C addersubtractor_0/fulladder_3/XOR_1/NAND_0/w_0_0# 0.06fF
C6 comparator_0/fourinputAND_1/fourinputNAND_0/a_76_n14# comparator_0/XNOR_1/out 0.23fF
C7 gnd twotofourdecoder_0/AND_2/not_0/in 0.04fF
C8 enableblock_2/enable1_1/AND_2/NAND_0/a_6_n14# enableblock_2/enable1_1/AND_2/not_0/in 0.12fF
C9 vdd addersubtractor_0/XOR_0/NAND_3/w_0_0# 0.05fF
C10 comparator_0/not_0/w_0_0# comparator_0/B3 0.06fF
C11 andblock_0/A1 andblock_0/AND_2/NAND_0/w_0_0# 0.06fF
C12 OR_0/in1 OR_0/NOR_0/w_0_0# 0.06fF
C13 comparator_0/A1 comparator_0/XNOR_2/XOR_0/NAND_1/w_0_0# 0.06fF
C14 comparator_0/XNOR_0/XOR_0/NAND_3/in1 comparator_0/XNOR_0/XOR_0/NAND_3/w_0_0# 0.06fF
C15 enableblock_2/enable1_1/AND_0/NAND_0/a_6_n14# enableblock_2/enable1_1/AND_0/not_0/in 0.12fF
C16 vdd enableblock_2/enable1_0/AND_0/not_0/in 0.29fF
C17 vdd twotofourdecoder_0/not_1/out 0.64fF
C18 vdd addersubtractor_0/XOR_1/NAND_3/in1 0.25fF
C19 addersubtractor_0/fulladder_1/OR_0/NOT_0/in addersubtractor_0/fulladder_1/OR_0/NOR_0/a_13_6# 0.04fF
C20 addersubtractor_0/fulladder_0/XOR_1/NAND_3/a_6_n14# gnd 0.57fF
C21 enableblock_2/En enableblock_2/enable1_0/AND_3/NAND_0/w_0_0# 0.06fF
C22 vdd addersubtractor_0/fulladder_0/XOR_1/NAND_3/w_32_0# 0.05fF
C23 S0 B1 0.16fF
C24 addersubtractor_0/fulladder_0/XOR_0/NAND_3/a_6_n14# gnd 0.57fF
C25 XOR_0/NAND_3/in1 XOR_0/NAND_3/w_0_0# 0.06fF
C26 gnd twotofourdecoder_0/AND_1/NAND_0/a_6_n14# 0.57fF
C27 addersubtractor_0/fulladder_0/XOR_1/NAND_0/a_6_n14# addersubtractor_0/fulladder_0/XOR_1/NAND_2/in1 0.12fF
C28 addersubtractor_0/fulladder_0/XOR_0/NAND_3/w_32_0# vdd 0.05fF
C29 comparator_0/A0 comparator_0/XNOR_3/XOR_0/NAND_1/w_0_0# 0.06fF
C30 comparator_0/XNOR_2/XOR_0/NAND_3/in1 comparator_0/XNOR_2/XOR_0/NAND_3/w_0_0# 0.06fF
C31 vdd twotofourdecoder_0/AND_0/not_0/w_0_0# 0.05fF
C32 enableblock_0/A_out3 S0 0.06fF
C33 addersubtractor_0/XOR_0/NAND_2/w_32_0# addersubtractor_0/XOR_0/NAND_3/in2 0.03fF
C34 enableblock_2/enable1_0/AND_3/NAND_0/w_32_0# enableblock_2/enable1_0/AND_3/not_0/in 0.03fF
C35 addersubtractor_0/fulladder_0/OR_0/in2 gnd 0.36fF
C36 gnd comparator_0/XNOR_3/out 0.10fF
C37 enableblock_1/enable1_1/AND_1/NAND_0/w_32_0# enableblock_1/enable1_1/AND_1/not_0/in 0.03fF
C38 addersubtractor_0/fulladder_1/OR_0/NOT_0/w_0_0# addersubtractor_0/fulladder_1/C 0.03fF
C39 comparator_0/threeinputAND_0/not_0/w_0_0# comparator_0/threeinputAND_0/not_0/in 0.06fF
C40 vdd Carry 0.25fF
C41 enableblock_0/enable1_0/AND_0/not_0/w_0_0# enableblock_0/enable1_0/AND_0/not_0/in 0.06fF
C42 enableblock_1/enable1_0/AND_3/not_0/in comparator_0/B2 0.02fF
C43 addersubtractor_0/fulladder_0/OR_0/in2 addersubtractor_0/fulladder_0/AND_0/not_0/in 0.02fF
C44 comparator_0/fourinputAND_1/fourinputNAND_0/w_63_0# comparator_0/fourinputAND_1/not_0/in 0.03fF
C45 vdd enableblock_2/enable1_1/AND_3/not_0/in 0.29fF
C46 addersubtractor_0/fulladder_1/XOR_1/NAND_0/a_6_n14# gnd 0.57fF
C47 addersubtractor_0/fulladder_0/XOR_1/NAND_2/in1 vdd 0.25fF
C48 vdd comparator_0/threeinputAND_0/not_0/in 1.58fF
C49 vdd enableblock_0/enable1_1/AND_3/NAND_0/w_32_0# 0.05fF
C50 vdd AND_0/not_0/w_0_0# 0.05fF
C51 addersubtractor_0/fulladder_2/XOR_1/NAND_3/w_0_0# adder2 0.03fF
C52 comparator_0/XNOR_3/XOR_0/NAND_3/in1 comparator_0/XNOR_3/XOR_0/NAND_3/w_0_0# 0.06fF
C53 enableblock_0/enable1_1/AND_3/NAND_0/w_32_0# B3 0.06fF
C54 addersubtractor_0/fulladder_2/OR_0/NOT_0/in addersubtractor_0/fulladder_2/OR_0/NOT_0/w_0_0# 0.06fF
C55 vdd addersubtractor_0/fulladder_2/XOR_1/NAND_3/in2 0.25fF
C56 gnd comparator_0/XNOR_1/XOR_0/NAND_2/in1 0.15fF
C57 addersubtractor_0/fulladder_2/XOR_1/NAND_2/in1 gnd 0.15fF
C58 vdd addersubtractor_0/fulladder_2/XOR_0/NAND_3/in2 0.25fF
C59 addersubtractor_0/fulladder_2/XOR_0/NAND_3/w_0_0# addersubtractor_0/fulladder_2/XOR_1/in2 0.03fF
C60 vdd comparator_0/XNOR_0/out 0.37fF
C61 gnd comparator_0/not_1/out 0.08fF
C62 vdd AND_0/NAND_0/w_32_0# 0.05fF
C63 enableblock_0/enable1_0/AND_3/not_0/w_0_0# enableblock_0/enable1_0/AND_3/not_0/in 0.06fF
C64 vdd enableblock_1/enable1_1/AND_2/NAND_0/w_0_0# 0.05fF
C65 gnd comparator_0/XNOR_0/XOR_0/NAND_0/a_6_n14# 0.57fF
C66 comparator_0/threeinputAND_0/threeinputNAND_0/a_6_n14# comparator_0/threeinputAND_0/not_0/in 0.11fF
C67 vdd enableblock_1/enable1_0/AND_0/NAND_0/w_0_0# 0.05fF
C68 enableblock_1/enable1_1/AND_0/not_0/w_0_0# enableblock_1/enable1_1/AND_0/not_0/in 0.06fF
C69 vdd addersubtractor_0/fulladder_1/XOR_1/NAND_0/w_0_0# 0.05fF
C70 OR_0/out OR_0/in1 0.06fF
C71 OR_0/NOT_0/in OR_0/NOT_0/w_0_0# 0.06fF
C72 vdd enableblock_0/enable1_0/AND_1/NAND_0/w_32_0# 0.05fF
C73 AND_2/in2 B1 0.06fF
C74 addersubtractor_0/fulladder_2/AND_1/NAND_0/w_32_0# addersubtractor_0/fulladder_2/XOR_1/in2 0.06fF
C75 addersubtractor_0/fulladder_1/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_1/XOR_1/NAND_0/w_0_0# 0.03fF
C76 B0 enableblock_2/enable1_1/AND_3/NAND_0/w_32_0# 0.06fF
C77 B2 enableblock_2/enable1_0/AND_3/NAND_0/w_32_0# 0.06fF
C78 gnd comparator_0/XNOR_2/XOR_0/NAND_0/a_6_n14# 0.57fF
C79 addersubtractor_0/XOR_2/NAND_3/in1 addersubtractor_0/XOR_2/NAND_1/w_0_0# 0.03fF
C80 vdd andblock_0/AND_0/not_0/w_0_0# 0.05fF
C81 gnd comparator_0/fourinputAND_0/fourinputNAND_0/a_6_n14# 0.47fF
C82 OR_0/out enableblock_0/enable1_1/AND_2/NAND_0/w_32_0# 0.06fF
C83 comparator_0/not_3/w_0_0# comparator_0/B0 0.06fF
C84 enableblock_1/enable1_1/AND_3/NAND_0/w_32_0# enableblock_1/enable1_1/AND_3/not_0/in 0.03fF
C85 gnd XOR_0/NAND_1/a_6_n14# 0.57fF
C86 comparator_0/fourinputOR_0/in4 comparator_0/XNOR_3/out 0.06fF
C87 gnd comparator_0/XNOR_3/XOR_0/NAND_0/a_6_n14# 0.57fF
C88 addersubtractor_0/XOR_3/out addersubtractor_0/XOR_3/NAND_3/a_6_n14# 0.12fF
C89 vdd addersubtractor_0/fulladder_3/OR_0/NOR_0/w_32_0# 0.03fF
C90 A0 A1 0.20fF
C91 vdd comparator_0/fiveinputAND_0/fiveinputNAND_0/w_63_0# 0.05fF
C92 enableblock_0/enable1_1/AND_1/NAND_0/a_6_n14# enableblock_0/enable1_1/AND_1/not_0/in 0.12fF
C93 vdd andblock_0/A1 0.20fF
C94 gnd enableblock_2/enable1_1/AND_0/NAND_0/a_6_n14# 0.57fF
C95 AND_0/not_0/w_0_0# XOR_0/in1 0.03fF
C96 gnd twotofourdecoder_0/not_0/out 0.42fF
C97 enableblock_2/enable1_1/AND_1/NAND_0/w_0_0# enableblock_2/enable1_1/AND_1/not_0/in 0.03fF
C98 addersubtractor_0/fulladder_0/XOR_1/in2 addersubtractor_0/fulladder_0/XOR_1/NAND_2/w_32_0# 0.06fF
C99 vdd comparator_0/XNOR_2/out 0.48fF
C100 gnd enableblock_1/enable1_0/AND_2/NAND_0/a_6_n14# 0.57fF
C101 comparator_0/XNOR_3/out comparator_0/XNOR_3/not_0/in 0.02fF
C102 comparator_0/fourinputAND_1/not_0/w_0_0# comparator_0/fourinputAND_1/not_0/in 0.06fF
C103 vdd enableblock_1/enable1_0/AND_1/not_0/w_0_0# 0.05fF
C104 comparator_0/fiveinputAND_0/not_0/in comparator_0/fiveinputAND_0/fiveinputNAND_0/w_133_0# 0.03fF
C105 addersubtractor_0/fulladder_0/XOR_0/NAND_0/a_6_n14# gnd 0.57fF
C106 comparator_0/fourinputAND_0/fourinputNAND_0/w_0_0# comparator_0/fourinputAND_0/not_0/in 0.03fF
C107 vdd enableblock_2/enable1_1/AND_0/NAND_0/w_32_0# 0.05fF
C108 addersubtractor_0/fulladder_2/AND_0/NAND_0/a_6_n14# gnd 0.57fF
C109 vdd addersubtractor_0/fulladder_1/OR_0/in2 0.07fF
C110 addersubtractor_0/XOR_0/NAND_3/in1 addersubtractor_0/XOR_0/NAND_3/w_0_0# 0.06fF
C111 addersubtractor_0/fulladder_1/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_1/XOR_1/NAND_1/a_6_n14# 0.12fF
C112 vdd enableblock_0/enable1_0/AND_3/NAND_0/w_0_0# 0.05fF
C113 addersubtractor_0/fulladder_0/AND_1/NAND_0/a_6_n14# addersubtractor_0/fulladder_0/AND_1/not_0/in 0.12fF
C114 enableblock_1/enable1_1/AND_1/not_0/in comparator_0/B1 0.02fF
C115 gnd enableblock_0/enable1_0/AND_0/not_0/in 0.04fF
C116 addersubtractor_0/fulladder_0/OR_0/NOR_0/a_13_6# addersubtractor_0/fulladder_0/OR_0/NOR_0/w_32_0# 0.03fF
C117 A0 S1 0.06fF
C118 vdd andblock_0/B1 0.20fF
C119 addersubtractor_0/fulladder_1/AND_1/not_0/in gnd 0.04fF
C120 addersubtractor_0/fulladder_1/XOR_0/NAND_3/in1 addersubtractor_0/fulladder_1/XOR_0/NAND_1/a_6_n14# 0.12fF
C121 comparator_0/XNOR_0/out comparator_0/fiveinputAND_0/fiveinputNAND_0/a_113_n14# 0.14fF
C122 gnd addersubtractor_0/fulladder_3/OR_0/in2 0.36fF
C123 vdd addersubtractor_0/fulladder_1/XOR_1/NAND_2/w_0_0# 0.05fF
C124 comparator_0/not_2/out comparator_0/XNOR_2/out 0.06fF
C125 addersubtractor_0/fulladder_2/XOR_1/NAND_1/w_32_0# addersubtractor_0/fulladder_2/XOR_1/NAND_3/in1 0.03fF
C126 addersubtractor_0/fulladder_1/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_1/XOR_1/NAND_2/w_0_0# 0.06fF
C127 addersubtractor_0/fulladder_3/AND_0/not_0/w_0_0# addersubtractor_0/fulladder_3/OR_0/in2 0.03fF
C128 addersubtractor_0/fulladder_1/XOR_1/in2 addersubtractor_0/fulladder_1/XOR_1/NAND_0/w_32_0# 0.06fF
C129 addersubtractor_0/fulladder_0/AND_0/NAND_0/w_32_0# addersubtractor_0/fulladder_0/AND_0/not_0/in 0.03fF
C130 vdd addersubtractor_0/fulladder_1/XOR_0/NAND_2/w_0_0# 0.05fF
C131 vdd enableblock_0/A_out1 0.32fF
C132 comparator_0/fourinputAND_0/fourinputNAND_0/a_45_n14# comparator_0/fourinputAND_0/fourinputNAND_0/a_76_n14# 0.04fF
C133 vdd addersubtractor_0/fulladder_2/XOR_0/NAND_2/in1 0.25fF
C134 addersubtractor_0/fulladder_2/XOR_1/NAND_2/w_0_0# addersubtractor_0/fulladder_2/XOR_1/NAND_3/in2 0.03fF
C135 gnd addersubtractor_0/fulladder_2/XOR_1/NAND_2/a_6_n14# 0.59fF
C136 addersubtractor_0/fulladder_2/XOR_0/NAND_1/w_32_0# addersubtractor_0/fulladder_2/XOR_0/NAND_3/in1 0.03fF
C137 vdd AND_2/in1 0.12fF
C138 A1 enableblock_2/enable1_1/AND_0/NAND_0/w_0_0# 0.06fF
C139 enableblock_2/enable1_0/AND_0/NAND_0/w_32_0# enableblock_2/En 0.06fF
C140 vdd addersubtractor_0/fulladder_2/XOR_1/NAND_2/w_32_0# 0.05fF
C141 vdd addersubtractor_0/fulladder_3/AND_0/not_0/in 0.29fF
C142 comparator_0/XNOR_3/XOR_0/NAND_2/in1 comparator_0/XNOR_3/XOR_0/NAND_0/a_6_n14# 0.12fF
C143 gnd enableblock_0/enable1_1/AND_3/not_0/in 0.04fF
C144 addersubtractor_0/fulladder_2/XOR_0/NAND_2/a_6_n14# gnd 0.59fF
C145 vdd addersubtractor_0/fulladder_1/OR_0/in1 0.12fF
C146 comparator_0/not_3/out comparator_0/fiveinputAND_0/fiveinputNAND_0/a_6_n14# 0.10fF
C147 vdd addersubtractor_0/fulladder_2/XOR_0/NAND_2/w_32_0# 0.05fF
C148 gnd enableblock_0/B_out1 1.65fF
C149 addersubtractor_0/fulladder_2/XOR_0/NAND_2/w_0_0# addersubtractor_0/fulladder_2/XOR_0/NAND_3/in2 0.03fF
C150 vdd addersubtractor_0/fulladder_2/XOR_0/NAND_0/w_0_0# 0.05fF
C151 enableblock_0/enable1_1/AND_3/NAND_0/a_6_n14# enableblock_0/enable1_1/AND_3/not_0/in 0.12fF
C152 vdd equal 0.09fF
C153 vdd addersubtractor_0/XOR_0/NAND_0/w_0_0# 0.05fF
C154 andblock_0/AND_2/not_0/in andblock_0/AND_2/NAND_0/w_0_0# 0.03fF
C155 addersubtractor_0/fulladder_2/OR_0/NOT_0/in addersubtractor_0/fulladder_2/C 0.02fF
C156 A1 A2 0.19fF
C157 gnd addersubtractor_0/XOR_1/NAND_2/in1 0.15fF
C158 addersubtractor_0/XOR_1/NAND_3/in1 addersubtractor_0/XOR_1/NAND_3/w_0_0# 0.06fF
C159 vdd comparator_0/fourinputOR_0/fourinputNOR_0/w_32_0# 0.03fF
C160 vdd addersubtractor_0/fulladder_3/OR_0/NOR_0/a_13_6# 0.21fF
C161 gnd addersubtractor_0/fulladder_3/OR_0/in1 0.30fF
C162 vdd andblock_0/AND_1/NAND_0/w_32_0# 0.05fF
C163 enableblock_1/enable1_0/AND_1/not_0/w_0_0# enableblock_1/enable1_0/AND_1/not_0/in 0.06fF
C164 vdd addersubtractor_0/XOR_3/out 0.32fF
C165 B2 enableblock_2/En 0.13fF
C166 vdd enableblock_1/enable1_1/AND_2/not_0/in 0.29fF
C167 comparator_0/threeinputAND_0/threeinputNAND_0/a_6_n14# comparator_0/threeinputAND_0/threeinputNAND_0/a_45_n14# 0.04fF
C168 gnd enableblock_2/enable1_0/AND_1/not_0/in 0.04fF
C169 vdd comparator_0/A3 0.32fF
C170 addersubtractor_0/fulladder_0/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_0/XOR_0/NAND_0/w_32_0# 0.03fF
C171 andblock_0/A3 andblock_0/AND_0/NAND_0/w_0_0# 0.06fF
C172 gnd addersubtractor_0/XOR_3/NAND_1/a_6_n14# 0.57fF
C173 vdd addersubtractor_0/XOR_3/NAND_1/w_32_0# 0.05fF
C174 comparator_0/fourinputOR_0/in3 comparator_0/fourinputAND_0/not_0/in 0.02fF
C175 vdd comparator_0/A1 0.20fF
C176 addersubtractor_0/XOR_3/NAND_3/w_32_0# addersubtractor_0/XOR_3/NAND_3/in2 0.06fF
C177 addersubtractor_0/fulladder_3/AND_1/NAND_0/w_32_0# addersubtractor_0/fulladder_3/AND_1/not_0/in 0.03fF
C178 comparator_0/XNOR_0/XOR_0/NAND_2/in1 comparator_0/XNOR_0/XOR_0/NAND_0/w_0_0# 0.03fF
C179 addersubtractor_0/XOR_0/NAND_3/in1 addersubtractor_0/XOR_0/NAND_1/a_6_n14# 0.12fF
C180 A2 S1 0.06fF
C181 vdd comparator_0/A0 0.26fF
C182 gnd addersubtractor_0/XOR_1/NAND_3/a_6_n14# 0.57fF
C183 vdd addersubtractor_0/XOR_1/NAND_3/w_32_0# 0.05fF
C184 A1 A3 0.19fF
C185 comparator_0/fiveinputAND_0/fiveinputNAND_0/w_32_0# comparator_0/A0 0.06fF
C186 addersubtractor_0/fulladder_2/AND_0/not_0/in addersubtractor_0/fulladder_2/AND_0/NAND_0/a_6_n14# 0.12fF
C187 comparator_0/fourinputOR_0/in4 comparator_0/fourinputOR_0/fourinputNOR_0/w_97_0# 0.06fF
C188 enableblock_0/A_out3 enableblock_0/enable1_0/AND_0/not_0/in 0.02fF
C189 vdd andblock_0/AND_0/NAND_0/w_0_0# 0.05fF
C190 addersubtractor_0/fulladder_0/AND_0/NAND_0/w_32_0# enableblock_0/A_out3 0.06fF
C191 andblock_0/B2 andblock_0/AND_1/NAND_0/w_32_0# 0.06fF
C192 vdd comparator_0/AND_0/NAND_0/w_0_0# 0.05fF
C193 vdd addersubtractor_0/XOR_3/NAND_0/w_32_0# 0.05fF
C194 addersubtractor_0/fulladder_1/AND_1/not_0/w_0_0# addersubtractor_0/fulladder_1/OR_0/in1 0.03fF
C195 vdd twotofourdecoder_0/AND_2/NAND_0/w_0_0# 0.05fF
C196 vdd enableblock_0/enable1_0/AND_3/not_0/in 0.29fF
C197 AND_0/not_0/in AND_0/not_0/w_0_0# 0.06fF
C198 addersubtractor_0/fulladder_0/AND_0/NAND_0/a_6_n14# addersubtractor_0/XOR_0/out 0.07fF
C199 vdd enableblock_1/enable1_0/AND_3/NAND_0/w_32_0# 0.05fF
C200 addersubtractor_0/fulladder_2/AND_0/NAND_0/a_6_n14# addersubtractor_0/XOR_2/out 0.07fF
C201 addersubtractor_0/fulladder_1/AND_1/NAND_0/w_0_0# addersubtractor_0/fulladder_1/AND_1/not_0/in 0.03fF
C202 comparator_0/fourinputAND_0/fourinputNAND_0/a_45_n14# comparator_0/A1 0.21fF
C203 gnd enableblock_2/enable1_1/AND_3/NAND_0/a_6_n14# 0.57fF
C204 vdd enableblock_2/enable1_1/AND_2/not_0/w_0_0# 0.05fF
C205 addersubtractor_0/fulladder_0/OR_0/NOT_0/in vdd 0.11fF
C206 addersubtractor_0/fulladder_0/C gnd 1.14fF
C207 gnd enableblock_0/B_out2 0.82fF
C208 A3 S1 0.06fF
C209 comparator_0/fourinputOR_0/fourinputNOR_0/a_45_6# comparator_0/fourinputOR_0/fourinputNOR_0/w_32_0# 0.03fF
C210 AND_0/not_0/in AND_0/NAND_0/w_32_0# 0.03fF
C211 addersubtractor_0/fulladder_2/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_2/XOR_0/NAND_2/w_0_0# 0.06fF
C212 vdd addersubtractor_0/fulladder_1/XOR_1/NAND_3/in1 0.25fF
C213 vdd enableblock_0/enable1_0/AND_0/NAND_0/w_32_0# 0.05fF
C214 addersubtractor_0/fulladder_2/OR_0/NOT_0/in gnd 0.60fF
C215 vdd addersubtractor_0/fulladder_1/XOR_0/NAND_3/in1 0.25fF
C216 vdd andblock_0/AND_2/not_0/in 0.29fF
C217 addersubtractor_0/XOR_1/NAND_0/w_0_0# enableblock_0/A_out0 0.06fF
C218 enableblock_0/enable1_1/AND_2/NAND_0/w_0_0# enableblock_0/enable1_1/AND_2/not_0/in 0.03fF
C219 enableblock_0/B_out3 addersubtractor_0/fulladder_2/XOR_0/NAND_0/w_0_0# 0.06fF
C220 comparator_0/XNOR_3/XOR_0/NAND_2/in1 comparator_0/XNOR_3/XOR_0/NAND_2/w_0_0# 0.06fF
C221 S0 twotofourdecoder_0/AND_0/NAND_0/a_6_n14# 0.11fF
C222 gnd addersubtractor_0/fulladder_3/XOR_1/NAND_3/in1 0.11fF
C223 vdd addersubtractor_0/fulladder_3/XOR_1/NAND_1/w_0_0# 0.05fF
C224 vdd comparator_0/AND_0/out 0.76fF
C225 gnd addersubtractor_0/fulladder_3/XOR_0/NAND_3/in1 0.11fF
C226 vdd addersubtractor_0/fulladder_3/XOR_0/NAND_1/w_0_0# 0.05fF
C227 comparator_0/XNOR_2/XOR_0/NAND_2/in1 comparator_0/XNOR_2/XOR_0/NAND_0/w_0_0# 0.03fF
C228 addersubtractor_0/fulladder_1/C addersubtractor_0/fulladder_2/XOR_1/in2 0.06fF
C229 gnd comparator_0/XNOR_1/XOR_0/NAND_3/in1 0.11fF
C230 addersubtractor_0/XOR_1/NAND_1/w_32_0# addersubtractor_0/XOR_1/NAND_2/in1 0.06fF
C231 vdd comparator_0/XNOR_1/XOR_0/NAND_1/w_0_0# 0.05fF
C232 vdd S0 0.51fF
C233 S0 B3 0.17fF
C234 vdd andblock_0/AND_2/NAND_0/w_32_0# 0.05fF
C235 twotofourdecoder_0/AND_2/not_0/w_0_0# twotofourdecoder_0/AND_2/not_0/in 0.06fF
C236 enableblock_2/En enableblock_2/enable1_1/AND_3/NAND_0/w_0_0# 0.06fF
C237 addersubtractor_0/XOR_0/NAND_3/w_32_0# addersubtractor_0/XOR_0/NAND_3/in2 0.06fF
C238 gnd comparator_0/XNOR_0/XOR_0/NAND_3/in1 0.11fF
C239 addersubtractor_0/fulladder_2/OR_0/NOT_0/in addersubtractor_0/fulladder_2/OR_0/NOR_0/w_32_0# 0.03fF
C240 AND_2/in2 enableblock_1/enable1_0/AND_1/NAND_0/w_0_0# 0.06fF
C241 addersubtractor_0/fulladder_0/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_0/XOR_0/NAND_1/w_32_0# 0.06fF
C242 gnd andblock_0/A2 0.36fF
C243 addersubtractor_0/XOR_3/out addersubtractor_0/fulladder_3/XOR_0/NAND_2/w_32_0# 0.06fF
C244 comparator_0/XNOR_1/XOR_0/NAND_2/in1 comparator_0/XNOR_1/XOR_0/NAND_1/w_32_0# 0.06fF
C245 gnd comparator_0/XNOR_2/XOR_0/NAND_3/in1 0.11fF
C246 twotofourdecoder_0/AND_3/NAND_0/a_6_n14# twotofourdecoder_0/not_1/out 0.07fF
C247 enableblock_1/enable1_0/AND_2/NAND_0/w_32_0# enableblock_1/enable1_0/AND_2/not_0/in 0.03fF
C248 addersubtractor_0/XOR_3/NAND_2/a_6_n14# addersubtractor_0/XOR_3/NAND_3/in2 0.12fF
C249 B0 B2 0.19fF
C250 andblock_0/A0 andblock_0/AND_3/NAND_0/a_6_n14# 0.02fF
C251 gnd comparator_0/XNOR_3/XOR_0/NAND_3/in1 0.11fF
C252 addersubtractor_0/fulladder_1/OR_0/in2 addersubtractor_0/fulladder_1/OR_0/NOT_0/in 0.26fF
C253 A0 A2 0.19fF
C254 OR_0/NOT_0/in OR_0/NOR_0/w_32_0# 0.03fF
C255 vdd enableblock_0/A_out2 0.29fF
C256 gnd A1 0.33fF
C257 vdd OR_0/NOT_0/in 0.11fF
C258 gnd enableblock_1/enable1_0/AND_0/not_0/in 0.04fF
C259 addersubtractor_0/fulladder_0/XOR_1/NAND_3/w_32_0# adder0 0.03fF
C260 gnd enableblock_1/enable1_1/AND_1/NAND_0/a_6_n14# 0.57fF
C261 addersubtractor_0/fulladder_0/XOR_0/NAND_3/w_32_0# addersubtractor_0/fulladder_0/XOR_1/in2 0.03fF
C262 vdd AND_2/in2 0.66fF
C263 vdd twotofourdecoder_0/AND_2/not_0/in 0.29fF
C264 AND_2/in2 B3 0.06fF
C265 addersubtractor_0/fulladder_1/AND_1/NAND_0/w_0_0# addersubtractor_0/fulladder_0/C 0.06fF
C266 comparator_0/fourinputAND_0/fourinputNAND_0/w_63_0# comparator_0/XNOR_1/out 0.06fF
C267 comparator_0/AND_0/NAND_0/w_32_0# comparator_0/A3 0.06fF
C268 gnd enableblock_1/enable1_0/AND_3/not_0/in 0.04fF
C269 gnd S1 0.78fF
C270 andblock_0/B0 enableblock_2/enable1_1/AND_3/not_0/in 0.02fF
C271 enableblock_1/enable1_1/AND_3/not_0/w_0_0# comparator_0/B0 0.03fF
C272 comparator_0/fourinputOR_0/not_0/in comparator_0/AND_0/out 0.67fF
C273 A0 A3 0.19fF
C274 vdd addersubtractor_0/fulladder_1/XOR_1/NAND_3/w_0_0# 0.05fF
C275 vdd XOR_0/NAND_3/in2 0.25fF
C276 comparator_0/fourinputAND_0/not_0/in comparator_0/XNOR_1/out 0.03fF
C277 addersubtractor_0/fulladder_1/XOR_1/in2 gnd 0.63fF
C278 vdd addersubtractor_0/fulladder_1/XOR_0/NAND_3/w_0_0# 0.05fF
C279 enableblock_2/enable1_0/AND_3/NAND_0/w_0_0# enableblock_2/enable1_0/AND_3/not_0/in 0.03fF
C280 OR_0/out B0 0.06fF
C281 and1 andblock_0/AND_2/not_0/w_0_0# 0.03fF
C282 gnd comparator_0/fourinputAND_1/not_0/in 0.01fF
C283 addersubtractor_0/fulladder_0/OR_0/in2 vdd 0.07fF
C284 enableblock_2/En twotofourdecoder_0/not_1/out 0.06fF
C285 vdd comparator_0/XNOR_3/out 0.36fF
C286 gnd enableblock_1/enable1_1/AND_2/NAND_0/a_6_n14# 0.57fF
C287 addersubtractor_0/fulladder_2/OR_0/NOT_0/in addersubtractor_0/fulladder_2/OR_0/NOR_0/a_13_6# 0.04fF
C288 vdd enableblock_1/enable1_1/AND_1/not_0/w_0_0# 0.05fF
C289 gnd addersubtractor_0/fulladder_2/XOR_1/NAND_3/a_6_n14# 0.57fF
C290 vdd addersubtractor_0/fulladder_2/XOR_1/NAND_3/w_32_0# 0.05fF
C291 enableblock_0/enable1_0/AND_2/NAND_0/a_6_n14# enableblock_0/enable1_0/AND_2/not_0/in 0.12fF
C292 gnd comparator_0/B2 0.22fF
C293 addersubtractor_0/fulladder_1/AND_1/NAND_0/w_32_0# vdd 0.05fF
C294 addersubtractor_0/fulladder_2/XOR_0/NAND_3/a_6_n14# gnd 0.57fF
C295 vdd addersubtractor_0/fulladder_2/XOR_0/NAND_3/w_32_0# 0.05fF
C296 addersubtractor_0/fulladder_1/XOR_1/NAND_0/a_6_n14# addersubtractor_0/fulladder_1/XOR_1/NAND_2/in1 0.12fF
C297 enableblock_2/En twotofourdecoder_0/AND_0/not_0/w_0_0# 0.03fF
C298 vdd enableblock_0/enable1_1/AND_3/NAND_0/w_0_0# 0.05fF
C299 addersubtractor_0/XOR_0/NAND_2/in1 addersubtractor_0/XOR_0/NAND_2/w_0_0# 0.06fF
C300 gnd AND_2/not_0/in 0.04fF
C301 enableblock_0/B_out3 S0 0.06fF
C302 addersubtractor_0/XOR_1/NAND_0/w_32_0# vdd 0.05fF
C303 addersubtractor_0/fulladder_2/OR_0/NOT_0/w_0_0# addersubtractor_0/fulladder_2/C 0.03fF
C304 A1 B1 0.23fF
C305 vdd comparator_0/XNOR_1/XOR_0/NAND_2/in1 0.25fF
C306 comparator_0/fourinputAND_1/fourinputNAND_0/a_45_n14# comparator_0/fourinputAND_1/fourinputNAND_0/a_76_n14# 0.04fF
C307 AND_2/not_0/w_0_0# AND_2/not_0/in 0.06fF
C308 gnd addersubtractor_0/fulladder_3/XOR_1/NAND_0/a_6_n14# 0.57fF
C309 vdd addersubtractor_0/fulladder_2/XOR_1/NAND_2/in1 0.25fF
C310 vdd comparator_0/not_1/out 0.07fF
C311 greater comparator_0/NOR_0/w_0_0# 0.06fF
C312 A2 enableblock_0/enable1_1/AND_0/NAND_0/a_6_n14# 0.07fF
C313 addersubtractor_0/fulladder_3/XOR_1/NAND_3/w_0_0# adder3 0.03fF
C314 addersubtractor_0/fulladder_3/OR_0/NOT_0/in addersubtractor_0/fulladder_3/OR_0/NOT_0/w_0_0# 0.06fF
C315 vdd comparator_0/fourinputAND_0/fourinputNAND_0/w_100_0# 0.05fF
C316 comparator_0/XNOR_1/XOR_0/NAND_2/in1 comparator_0/XNOR_1/XOR_0/NAND_0/a_6_n14# 0.12fF
C317 vdd enableblock_2/enable1_0/AND_1/NAND_0/w_0_0# 0.05fF
C318 gnd addersubtractor_0/XOR_3/NAND_3/in1 0.11fF
C319 addersubtractor_0/XOR_0/out addersubtractor_0/XOR_0/NAND_3/w_32_0# 0.03fF
C320 gnd comparator_0/not_3/out 0.35fF
C321 twotofourdecoder_0/not_1/out twotofourdecoder_0/not_1/w_0_0# 0.03fF
C322 twotofourdecoder_0/AND_3/NAND_0/w_32_0# twotofourdecoder_0/AND_3/not_0/in 0.03fF
C323 S0 addersubtractor_0/XOR_2/NAND_2/w_32_0# 0.06fF
C324 gnd and1 0.08fF
C325 AND_2/NAND_0/w_0_0# AND_2/in1 0.06fF
C326 addersubtractor_0/fulladder_0/XOR_1/NAND_2/w_32_0# addersubtractor_0/fulladder_0/XOR_1/NAND_3/in2 0.03fF
C327 addersubtractor_0/fulladder_3/XOR_0/NAND_3/w_0_0# addersubtractor_0/fulladder_3/XOR_1/in2 0.03fF
C328 comparator_0/fourinputOR_0/in4 comparator_0/fiveinputAND_0/not_0/w_0_0# 0.03fF
C329 comparator_0/fourinputAND_1/fourinputNAND_0/w_100_0# comparator_0/XNOR_2/out 0.06fF
C330 gnd comparator_0/not_0/out 0.08fF
C331 enableblock_1/enable1_1/AND_3/NAND_0/w_0_0# enableblock_1/enable1_1/AND_3/not_0/in 0.03fF
C332 B1 S1 0.06fF
C333 andblock_0/AND_3/not_0/in andblock_0/AND_3/NAND_0/w_0_0# 0.03fF
C334 comparator_0/not_1/out comparator_0/threeinputAND_0/threeinputNAND_0/a_6_n14# 0.02fF
C335 gnd enableblock_0/enable1_0/AND_3/NAND_0/a_6_n14# 0.57fF
C336 vdd enableblock_0/enable1_0/AND_2/not_0/w_0_0# 0.05fF
C337 gnd comparator_0/fiveinputAND_0/fiveinputNAND_0/a_6_n14# 0.35fF
C338 vdd addersubtractor_0/fulladder_3/XOR_1/NAND_0/w_0_0# 0.05fF
C339 A2 A3 0.19fF
C340 gnd XOR_0/NAND_0/a_6_n14# 0.57fF
C341 comparator_0/fourinputAND_0/not_0/in comparator_0/XNOR_0/out 0.01fF
C342 addersubtractor_0/XOR_1/NAND_2/in1 addersubtractor_0/XOR_1/NAND_2/w_0_0# 0.06fF
C343 addersubtractor_0/fulladder_2/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_2/XOR_1/NAND_0/w_0_0# 0.03fF
C344 addersubtractor_0/fulladder_0/XOR_0/NAND_2/w_32_0# addersubtractor_0/fulladder_0/XOR_0/NAND_3/in2 0.03fF
C345 vdd andblock_0/AND_3/NAND_0/w_0_0# 0.05fF
C346 comparator_0/XNOR_0/XOR_0/NAND_1/w_0_0# comparator_0/XNOR_0/XOR_0/NAND_3/in1 0.03fF
C347 enableblock_2/enable1_1/AND_0/NAND_0/w_0_0# enableblock_2/enable1_1/AND_0/not_0/in 0.03fF
C348 addersubtractor_0/fulladder_3/AND_1/NAND_0/w_32_0# addersubtractor_0/fulladder_3/XOR_1/in2 0.06fF
C349 gnd andblock_0/AND_3/NAND_0/a_6_n14# 0.57fF
C350 comparator_0/XNOR_1/XOR_0/NAND_3/w_0_0# comparator_0/XNOR_1/not_0/in 0.03fF
C351 comparator_0/fiveinputAND_0/not_0/in comparator_0/fiveinputAND_0/fiveinputNAND_0/w_63_0# 0.03fF
C352 enableblock_2/enable1_1/AND_2/not_0/w_0_0# enableblock_2/enable1_1/AND_2/not_0/in 0.06fF
C353 comparator_0/A2 comparator_0/B3 2.23fF
C354 vdd comparator_0/fourinputAND_1/fourinputNAND_0/w_32_0# 0.05fF
C355 vdd andblock_0/AND_1/not_0/w_0_0# 0.05fF
C356 vdd twotofourdecoder_0/not_0/out 0.13fF
C357 addersubtractor_0/fulladder_0/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_0/XOR_1/NAND_0/w_32_0# 0.03fF
C358 vdd andblock_0/AND_1/NAND_0/w_0_0# 0.05fF
C359 enableblock_1/enable1_0/AND_0/not_0/w_0_0# comparator_0/A3 0.03fF
C360 gnd enableblock_2/enable1_1/AND_1/not_0/in 0.04fF
C361 enableblock_2/enable1_0/AND_0/NAND_0/a_6_n14# enableblock_2/enable1_0/AND_0/not_0/in 0.12fF
C362 addersubtractor_0/XOR_0/out gnd 0.56fF
C363 comparator_0/not_2/out comparator_0/fourinputAND_0/fourinputNAND_0/a_6_n14# 0.02fF
C364 comparator_0/fiveinputAND_0/not_0/in comparator_0/XNOR_2/out 0.16fF
C365 enableblock_2/enable1_0/AND_0/not_0/w_0_0# andblock_0/A3 0.03fF
C366 comparator_0/XNOR_2/XOR_0/NAND_1/w_0_0# comparator_0/XNOR_2/XOR_0/NAND_3/in1 0.03fF
C367 vdd addersubtractor_0/fulladder_1/AND_0/NAND_0/w_32_0# 0.05fF
C368 gnd XOR_0/NAND_2/a_6_n14# 0.59fF
C369 comparator_0/XNOR_0/XOR_0/NAND_3/w_0_0# comparator_0/XNOR_0/not_0/in 0.03fF
C370 addersubtractor_0/fulladder_1/XOR_1/in2 addersubtractor_0/fulladder_1/XOR_1/NAND_2/w_32_0# 0.06fF
C371 vdd XOR_0/NAND_2/w_32_0# 0.05fF
C372 enableblock_0/B_out2 enableblock_0/enable1_1/AND_1/not_0/in 0.02fF
C373 addersubtractor_0/fulladder_0/OR_0/NOT_0/w_0_0# vdd 0.05fF
C374 vdd enableblock_0/enable1_0/AND_0/not_0/in 0.29fF
C375 gnd A0 0.23fF
C376 OR_0/NOR_0/a_13_6# OR_0/NOR_0/w_32_0# 0.03fF
C377 comparator_0/fourinputAND_0/fourinputNAND_0/a_6_n14# comparator_0/fourinputAND_0/fourinputNAND_0/a_45_n14# 0.04fF
C378 addersubtractor_0/fulladder_2/XOR_0/NAND_0/a_6_n14# gnd 0.57fF
C379 vdd addersubtractor_0/fulladder_2/AND_1/not_0/w_0_0# 0.05fF
C380 vdd addersubtractor_0/fulladder_1/AND_1/not_0/in 0.29fF
C381 addersubtractor_0/fulladder_0/AND_0/NAND_0/a_6_n14# gnd 0.57fF
C382 vdd OR_0/NOR_0/a_13_6# 0.21fF
C383 comparator_0/fourinputOR_0/in4 comparator_0/not_3/out 0.04fF
C384 enableblock_2/En enableblock_2/enable1_1/AND_0/NAND_0/w_32_0# 0.06fF
C385 vdd addersubtractor_0/fulladder_3/OR_0/in2 0.07fF
C386 addersubtractor_0/fulladder_0/AND_0/NAND_0/w_32_0# vdd 0.05fF
C387 gnd addersubtractor_0/XOR_0/NAND_0/a_6_n14# 0.57fF
C388 addersubtractor_0/fulladder_2/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_2/XOR_1/NAND_1/a_6_n14# 0.12fF
C389 comparator_0/NOR_0/w_0_0# comparator_0/NOR_0/a_13_6# 0.03fF
C390 comparator_0/XNOR_3/XOR_0/NAND_1/w_0_0# comparator_0/XNOR_3/XOR_0/NAND_3/in1 0.03fF
C391 comparator_0/XNOR_1/XOR_0/NAND_0/w_32_0# comparator_0/XNOR_1/XOR_0/NAND_2/in1 0.03fF
C392 addersubtractor_0/fulladder_0/AND_0/NAND_0/a_6_n14# addersubtractor_0/fulladder_0/AND_0/not_0/in 0.12fF
C393 comparator_0/XNOR_2/XOR_0/NAND_3/w_0_0# comparator_0/XNOR_2/not_0/in 0.03fF
C394 enableblock_0/enable1_0/AND_1/NAND_0/w_0_0# enableblock_0/enable1_0/AND_1/not_0/in 0.03fF
C395 vdd addersubtractor_0/fulladder_1/OR_0/NOR_0/w_0_0# 0.05fF
C396 vdd comparator_0/fourinputOR_0/fourinputNOR_0/a_13_6# 0.21fF
C397 gnd enableblock_2/enable1_0/AND_1/NAND_0/a_6_n14# 0.57fF
C398 addersubtractor_0/fulladder_1/OR_0/NOR_0/a_13_6# addersubtractor_0/fulladder_1/OR_0/NOR_0/w_32_0# 0.03fF
C399 vdd enableblock_2/enable1_0/AND_0/not_0/w_0_0# 0.05fF
C400 gnd addersubtractor_0/fulladder_3/AND_1/not_0/in 0.04fF
C401 comparator_0/NOR_0/w_32_0# comparator_0/NOR_0/a_13_6# 0.03fF
C402 vdd addersubtractor_0/XOR_0/NAND_1/w_0_0# 0.05fF
C403 addersubtractor_0/fulladder_2/XOR_0/NAND_3/in1 addersubtractor_0/fulladder_2/XOR_0/NAND_1/a_6_n14# 0.12fF
C404 OR_0/out OR_0/in2 0.76fF
C405 vdd addersubtractor_0/fulladder_3/XOR_1/NAND_2/w_0_0# 0.05fF
C406 addersubtractor_0/fulladder_3/XOR_1/NAND_1/w_32_0# addersubtractor_0/fulladder_3/XOR_1/NAND_3/in1 0.03fF
C407 addersubtractor_0/fulladder_2/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_2/XOR_1/NAND_2/w_0_0# 0.06fF
C408 addersubtractor_0/fulladder_2/XOR_1/in2 addersubtractor_0/fulladder_2/XOR_1/NAND_0/w_32_0# 0.06fF
C409 vdd comparator_0/fourinputOR_0/fourinputNOR_0/w_97_0# 0.03fF
C410 vdd enableblock_0/enable1_1/AND_3/not_0/in 0.29fF
C411 vdd addersubtractor_0/fulladder_3/XOR_0/NAND_2/w_0_0# 0.05fF
C412 comparator_0/XNOR_3/XOR_0/NAND_3/w_0_0# comparator_0/XNOR_3/not_0/in 0.03fF
C413 vdd enableblock_1/enable1_1/AND_3/NAND_0/w_32_0# 0.05fF
C414 vdd enableblock_0/B_out1 0.29fF
C415 vdd comparator_0/XNOR_1/XOR_0/NAND_2/w_0_0# 0.05fF
C416 vdd addersubtractor_0/XOR_1/NAND_2/in1 0.25fF
C417 addersubtractor_0/fulladder_3/XOR_1/NAND_2/w_0_0# addersubtractor_0/fulladder_3/XOR_1/NAND_3/in2 0.03fF
C418 addersubtractor_0/fulladder_3/XOR_0/NAND_1/w_32_0# addersubtractor_0/fulladder_3/XOR_0/NAND_3/in1 0.03fF
C419 enableblock_2/enable1_1/AND_1/NAND_0/w_32_0# enableblock_2/enable1_1/AND_1/not_0/in 0.03fF
C420 gnd addersubtractor_0/XOR_3/NAND_2/in1 0.15fF
C421 vdd addersubtractor_0/XOR_2/NAND_2/w_0_0# 0.05fF
C422 comparator_0/fiveinputAND_0/fiveinputNAND_0/a_76_n14# comparator_0/fiveinputAND_0/fiveinputNAND_0/a_113_n14# 0.04fF
C423 twotofourdecoder_0/AND_0/not_0/w_0_0# twotofourdecoder_0/AND_0/not_0/in 0.06fF
C424 vdd addersubtractor_0/fulladder_3/OR_0/in1 0.12fF
C425 comparator_0/not_2/w_0_0# comparator_0/B1 0.06fF
C426 vdd comparator_0/XNOR_0/XOR_0/NAND_2/w_0_0# 0.05fF
C427 addersubtractor_0/XOR_2/out addersubtractor_0/XOR_2/NAND_3/w_0_0# 0.03fF
C428 addersubtractor_0/fulladder_3/XOR_0/NAND_2/w_0_0# addersubtractor_0/fulladder_3/XOR_0/NAND_3/in2 0.03fF
C429 comparator_0/XNOR_1/XOR_0/NAND_1/w_32_0# comparator_0/XNOR_1/XOR_0/NAND_3/in1 0.03fF
C430 enableblock_2/enable1_1/AND_1/not_0/w_0_0# andblock_0/B1 0.03fF
C431 addersubtractor_0/fulladder_0/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_0/XOR_0/NAND_0/w_0_0# 0.03fF
C432 vdd enableblock_2/enable1_0/AND_1/not_0/in 0.29fF
C433 vdd comparator_0/XNOR_2/XOR_0/NAND_2/w_0_0# 0.05fF
C434 AND_2/in2 OR_0/in1 0.13fF
C435 enableblock_0/A_out1 enableblock_0/enable1_0/AND_2/not_0/in 0.02fF
C436 comparator_0/XNOR_1/XOR_0/NAND_2/w_0_0# comparator_0/XNOR_1/XOR_0/NAND_3/in2 0.03fF
C437 enableblock_0/A_out3 addersubtractor_0/XOR_0/out 0.11fF
C438 gnd lesser 0.41fF
C439 gnd twotofourdecoder_0/AND_2/NAND_0/a_6_n14# 0.57fF
C440 vdd twotofourdecoder_0/AND_1/not_0/w_0_0# 0.05fF
C441 twotofourdecoder_0/AND_1/NAND_0/w_32_0# twotofourdecoder_0/not_0/out 0.06fF
C442 gnd A2 0.32fF
C443 vdd comparator_0/XNOR_3/XOR_0/NAND_2/w_0_0# 0.05fF
C444 addersubtractor_0/fulladder_1/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_1/XOR_0/NAND_0/w_32_0# 0.03fF
C445 addersubtractor_0/fulladder_1/AND_1/not_0/w_0_0# addersubtractor_0/fulladder_1/AND_1/not_0/in 0.06fF
C446 addersubtractor_0/fulladder_0/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_0/XOR_1/NAND_1/w_32_0# 0.06fF
C447 enableblock_1/enable1_0/AND_3/NAND_0/a_6_n14# enableblock_1/enable1_0/AND_3/not_0/in 0.12fF
C448 A0 B1 3.14fF
C449 addersubtractor_0/XOR_2/NAND_2/w_0_0# addersubtractor_0/XOR_2/NAND_3/in2 0.03fF
C450 gnd addersubtractor_0/XOR_2/NAND_0/a_6_n14# 0.57fF
C451 enableblock_2/enable1_1/AND_0/not_0/w_0_0# enableblock_2/enable1_1/AND_0/not_0/in 0.06fF
C452 comparator_0/fourinputOR_0/fourinputNOR_0/a_45_6# comparator_0/fourinputOR_0/fourinputNOR_0/a_13_6# 0.04fF
C453 gnd enableblock_0/enable1_1/AND_0/NAND_0/a_6_n14# 0.57fF
C454 comparator_0/XNOR_0/XOR_0/NAND_2/w_0_0# comparator_0/XNOR_0/XOR_0/NAND_3/in2 0.03fF
C455 vdd twotofourdecoder_0/AND_0/NAND_0/w_0_0# 0.05fF
C456 AND_2/in2 enableblock_1/enable1_1/AND_1/NAND_0/w_0_0# 0.06fF
C457 enableblock_2/enable1_1/AND_3/NAND_0/w_32_0# enableblock_2/enable1_1/AND_3/not_0/in 0.03fF
C458 gnd andblock_0/A0 0.53fF
C459 enableblock_0/enable1_0/AND_1/NAND_0/w_32_0# B0 0.06fF
C460 andblock_0/A2 enableblock_2/enable1_0/AND_2/not_0/in 0.02fF
C461 A3 enableblock_2/enable1_0/AND_0/NAND_0/w_0_0# 0.06fF
C462 enableblock_0/enable1_0/AND_0/not_0/in enableblock_0/enable1_0/AND_0/NAND_0/w_0_0# 0.03fF
C463 vdd enableblock_0/enable1_1/AND_0/NAND_0/w_32_0# 0.05fF
C464 AND_2/NAND_0/a_6_n14# AND_2/not_0/in 0.12fF
C465 addersubtractor_0/fulladder_3/AND_0/not_0/in addersubtractor_0/fulladder_3/AND_0/NAND_0/a_6_n14# 0.12fF
C466 andblock_0/AND_1/not_0/in andblock_0/AND_1/NAND_0/w_32_0# 0.03fF
C467 vdd enableblock_1/enable1_0/AND_3/NAND_0/w_0_0# 0.05fF
C468 enableblock_1/enable1_0/AND_2/not_0/in comparator_0/A2 0.02fF
C469 comparator_0/XNOR_2/XOR_0/NAND_2/w_0_0# comparator_0/XNOR_2/XOR_0/NAND_3/in2 0.03fF
C470 vdd addersubtractor_0/fulladder_0/C 0.18fF
C471 comparator_0/fourinputOR_0/not_0/in comparator_0/fourinputOR_0/fourinputNOR_0/w_97_0# 0.03fF
C472 vdd enableblock_0/B_out2 0.20fF
C473 gnd A3 0.32fF
C474 addersubtractor_0/fulladder_2/AND_1/not_0/w_0_0# addersubtractor_0/fulladder_2/OR_0/in1 0.03fF
C475 gnd comparator_0/AND_0/not_0/in 0.04fF
C476 addersubtractor_0/fulladder_3/AND_0/NAND_0/a_6_n14# addersubtractor_0/XOR_3/out 0.07fF
C477 addersubtractor_0/fulladder_0/XOR_1/in2 S0 0.06fF
C478 gnd andblock_0/AND_0/not_0/in 0.04fF
C479 comparator_0/XNOR_3/XOR_0/NAND_2/in1 comparator_0/XNOR_3/XOR_0/NAND_0/w_32_0# 0.03fF
C480 comparator_0/fiveinputAND_0/fiveinputNAND_0/a_45_n14# comparator_0/A0 0.14fF
C481 enableblock_0/enable1_1/AND_0/NAND_0/w_32_0# enableblock_0/enable1_1/AND_0/not_0/in 0.03fF
C482 vdd addersubtractor_0/fulladder_2/OR_0/NOT_0/in 0.11fF
C483 gnd addersubtractor_0/fulladder_2/C 1.20fF
C484 gnd enableblock_2/enable1_1/AND_0/not_0/in 0.04fF
C485 enableblock_0/enable1_1/AND_3/not_0/w_0_0# enableblock_0/enable1_1/AND_3/not_0/in 0.06fF
C486 comparator_0/XNOR_3/XOR_0/NAND_2/w_0_0# comparator_0/XNOR_3/XOR_0/NAND_3/in2 0.03fF
C487 addersubtractor_0/XOR_0/NAND_3/in1 addersubtractor_0/XOR_0/NAND_1/w_0_0# 0.03fF
C488 vdd addersubtractor_0/fulladder_3/XOR_1/NAND_3/in1 0.25fF
C489 addersubtractor_0/fulladder_3/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_3/XOR_0/NAND_2/w_0_0# 0.06fF
C490 addersubtractor_0/XOR_0/NAND_2/in1 addersubtractor_0/XOR_0/NAND_0/w_32_0# 0.03fF
C491 gnd enableblock_1/enable1_1/AND_3/not_0/in 0.04fF
C492 vdd addersubtractor_0/fulladder_3/XOR_0/NAND_3/in1 0.25fF
C493 addersubtractor_0/fulladder_0/AND_1/NAND_0/w_0_0# S0 0.06fF
C494 and3 andblock_0/AND_0/not_0/in 0.02fF
C495 comparator_0/not_1/w_0_0# comparator_0/not_1/out 0.03fF
C496 B1 A2 0.23fF
C497 vdd addersubtractor_0/XOR_3/NAND_3/in2 0.25fF
C498 vdd comparator_0/XNOR_1/XOR_0/NAND_3/in1 0.25fF
C499 enableblock_0/B_out1 addersubtractor_0/fulladder_3/XOR_0/NAND_0/w_0_0# 0.06fF
C500 addersubtractor_0/XOR_3/NAND_0/w_0_0# enableblock_0/B_out0 0.06fF
C501 vdd comparator_0/XNOR_0/XOR_0/NAND_3/in1 0.25fF
C502 addersubtractor_0/fulladder_2/C addersubtractor_0/fulladder_3/XOR_1/in2 0.06fF
C503 enableblock_0/A_out3 addersubtractor_0/fulladder_0/XOR_0/NAND_1/w_0_0# 0.06fF
C504 vdd andblock_0/A2 0.20fF
C505 OR_0/out B2 0.06fF
C506 S0 enableblock_2/En 0.75fF
C507 gnd enableblock_0/enable1_0/AND_1/not_0/in 0.04fF
C508 enableblock_1/enable1_1/AND_0/NAND_0/a_6_n14# A1 0.07fF
C509 vdd comparator_0/XNOR_2/XOR_0/NAND_3/in1 0.25fF
C510 enableblock_1/enable1_0/AND_2/NAND_0/w_0_0# enableblock_1/enable1_0/AND_2/not_0/in 0.03fF
C511 vdd addersubtractor_0/XOR_2/NAND_0/w_0_0# 0.05fF
C512 addersubtractor_0/fulladder_0/XOR_1/NAND_3/w_32_0# addersubtractor_0/fulladder_0/XOR_1/NAND_3/in2 0.06fF
C513 comparator_0/fourinputOR_0/in2 comparator_0/XNOR_1/out 0.06fF
C514 addersubtractor_0/fulladder_3/OR_0/NOT_0/in addersubtractor_0/fulladder_3/OR_0/NOR_0/w_32_0# 0.03fF
C515 vdd comparator_0/XNOR_3/XOR_0/NAND_3/in1 0.25fF
C516 enableblock_2/enable1_0/AND_1/not_0/w_0_0# enableblock_2/enable1_0/AND_1/not_0/in 0.06fF
C517 addersubtractor_0/fulladder_1/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_1/XOR_0/NAND_1/w_32_0# 0.06fF
C518 OR_0/in1 XOR_0/NAND_2/w_32_0# 0.06fF
C519 addersubtractor_0/fulladder_0/XOR_0/NAND_3/w_32_0# addersubtractor_0/fulladder_0/XOR_0/NAND_3/in2 0.06fF
C520 B1 A3 0.19fF
C521 A1 B3 0.19fF
C522 vdd enableblock_1/enable1_0/AND_0/not_0/in 0.29fF
C523 adder0 addersubtractor_0/fulladder_0/XOR_1/NAND_3/a_6_n14# 0.12fF
C524 vdd addersubtractor_0/XOR_0/NAND_3/in2 0.25fF
C525 vdd twotofourdecoder_0/AND_3/NAND_0/w_32_0# 0.05fF
C526 XOR_0/NAND_3/w_0_0# Carry 0.03fF
C527 addersubtractor_0/fulladder_2/OR_0/in2 addersubtractor_0/fulladder_2/OR_0/NOT_0/in 0.26fF
C528 comparator_0/XNOR_2/out comparator_0/XNOR_2/not_0/w_0_0# 0.03fF
C529 enableblock_1/enable1_0/AND_0/NAND_0/a_6_n14# enableblock_1/enable1_0/AND_0/not_0/in 0.12fF
C530 addersubtractor_0/fulladder_0/XOR_1/in2 addersubtractor_0/fulladder_0/XOR_0/NAND_3/a_6_n14# 0.12fF
C531 enableblock_1/enable1_1/AND_0/not_0/in comparator_0/A1 0.02fF
C532 addersubtractor_0/fulladder_1/AND_0/not_0/w_0_0# vdd 0.05fF
C533 vdd enableblock_2/enable1_1/AND_1/NAND_0/w_0_0# 0.05fF
C534 addersubtractor_0/fulladder_1/XOR_1/NAND_3/w_32_0# adder1 0.03fF
C535 andblock_0/AND_2/NAND_0/a_6_n14# andblock_0/AND_2/not_0/in 0.12fF
C536 enableblock_0/B_out3 enableblock_0/B_out2 0.78fF
C537 gnd XOR_0/NAND_3/a_6_n14# 0.57fF
C538 vdd XOR_0/NAND_3/w_32_0# 0.05fF
C539 enableblock_0/A_out3 enableblock_0/enable1_0/AND_0/not_0/w_0_0# 0.03fF
C540 vdd enableblock_1/enable1_0/AND_3/not_0/in 0.29fF
C541 vdd S1 0.13fF
C542 comparator_0/XNOR_0/XOR_0/NAND_1/w_32_0# comparator_0/XNOR_0/XOR_0/NAND_3/in1 0.03fF
C543 gnd enableblock_0/enable1_1/AND_3/NAND_0/a_6_n14# 0.57fF
C544 addersubtractor_0/fulladder_1/XOR_0/NAND_3/w_32_0# addersubtractor_0/fulladder_1/XOR_1/in2 0.03fF
C545 B3 S1 0.06fF
C546 S0 twotofourdecoder_0/not_0/w_0_0# 0.06fF
C547 vdd enableblock_0/enable1_1/AND_2/not_0/w_0_0# 0.05fF
C548 vdd addersubtractor_0/XOR_1/NAND_1/w_0_0# 0.05fF
C549 addersubtractor_0/fulladder_0/AND_0/not_0/in gnd 0.04fF
C550 vdd comparator_0/fourinputAND_1/fourinputNAND_0/w_63_0# 0.05fF
C551 comparator_0/threeinputAND_0/not_0/in comparator_0/fourinputOR_0/in2 0.02fF
C552 A2 enableblock_2/enable1_0/AND_2/NAND_0/w_0_0# 0.06fF
C553 vdd adder1 0.25fF
C554 addersubtractor_0/fulladder_0/OR_0/NOR_0/w_32_0# vdd 0.03fF
C555 vdd addersubtractor_0/fulladder_1/XOR_1/in2 0.47fF
C556 gnd and3 0.08fF
C557 vdd comparator_0/fiveinputAND_0/not_0/w_0_0# 0.05fF
C558 AND_2/NAND_0/w_32_0# AND_2/in2 0.06fF
C559 comparator_0/B1 comparator_0/XNOR_1/out 0.07fF
C560 comparator_0/XNOR_2/XOR_0/NAND_1/w_32_0# comparator_0/XNOR_2/XOR_0/NAND_3/in1 0.03fF
C561 enableblock_1/enable1_1/AND_1/not_0/w_0_0# enableblock_1/enable1_1/AND_1/not_0/in 0.06fF
C562 vdd comparator_0/fourinputAND_1/not_0/in 1.27fF
C563 enableblock_1/enable1_1/AND_0/not_0/w_0_0# comparator_0/A1 0.03fF
C564 gnd addersubtractor_0/XOR_3/NAND_2/a_6_n14# 0.59fF
C565 addersubtractor_0/XOR_0/NAND_2/a_6_n14# addersubtractor_0/XOR_0/NAND_3/in2 0.12fF
C566 andblock_0/AND_1/not_0/w_0_0# and2 0.03fF
C567 comparator_0/threeinputAND_0/threeinputNAND_0/w_0_0# comparator_0/threeinputAND_0/not_0/in 0.03fF
C568 vdd addersubtractor_0/XOR_3/NAND_2/w_32_0# 0.05fF
C569 vdd addersubtractor_0/fulladder_3/XOR_1/NAND_3/w_0_0# 0.05fF
C570 comparator_0/fourinputAND_1/fourinputNAND_0/a_6_n14# comparator_0/fourinputAND_1/fourinputNAND_0/a_45_n14# 0.04fF
C571 vdd comparator_0/B2 0.30fF
C572 addersubtractor_0/fulladder_2/AND_1/NAND_0/a_6_n14# gnd 0.57fF
C573 comparator_0/B0 comparator_0/XNOR_1/out 0.07fF
C574 vdd addersubtractor_0/fulladder_3/XOR_0/NAND_3/w_0_0# 0.05fF
C575 gnd addersubtractor_0/fulladder_3/XOR_1/in2 0.63fF
C576 comparator_0/XNOR_0/out comparator_0/A2 0.06fF
C577 vdd comparator_0/threeinputAND_0/threeinputNAND_0/w_32_0# 0.05fF
C578 enableblock_0/A_out0 enableblock_0/enable1_0/AND_3/not_0/in 0.02fF
C579 AND_2/in2 enableblock_1/enable1_0/AND_2/NAND_0/w_32_0# 0.06fF
C580 vdd AND_2/not_0/in 0.29fF
C581 gnd comparator_0/XNOR_1/not_0/in 0.03fF
C582 vdd addersubtractor_0/XOR_0/NAND_2/w_32_0# 0.05fF
C583 addersubtractor_0/fulladder_3/OR_0/NOT_0/in addersubtractor_0/fulladder_3/OR_0/NOR_0/a_13_6# 0.04fF
C584 addersubtractor_0/fulladder_0/XOR_1/NAND_1/w_0_0# addersubtractor_0/fulladder_0/XOR_1/NAND_3/in1 0.03fF
C585 comparator_0/XNOR_3/XOR_0/NAND_1/w_32_0# comparator_0/XNOR_3/XOR_0/NAND_3/in1 0.03fF
C586 vdd comparator_0/XNOR_1/XOR_0/NAND_3/w_0_0# 0.05fF
C587 comparator_0/threeinputAND_0/threeinputNAND_0/w_63_0# comparator_0/threeinputAND_0/not_0/in 0.03fF
C588 vdd comparator_0/fourinputAND_0/fourinputNAND_0/w_32_0# 0.05fF
C589 andblock_0/B3 andblock_0/AND_0/NAND_0/w_32_0# 0.06fF
C590 enableblock_2/enable1_0/AND_0/NAND_0/w_32_0# enableblock_2/enable1_0/AND_0/not_0/in 0.03fF
C591 vdd addersubtractor_0/XOR_2/NAND_3/w_0_0# 0.05fF
C592 addersubtractor_0/XOR_1/NAND_1/a_6_n14# addersubtractor_0/XOR_1/NAND_3/in1 0.12fF
C593 vdd addersubtractor_0/fulladder_3/AND_1/NAND_0/w_32_0# 0.05fF
C594 gnd comparator_0/XNOR_0/not_0/in 0.03fF
C595 gnd comparator_0/fourinputOR_0/in4 0.21fF
C596 addersubtractor_0/fulladder_2/XOR_1/NAND_0/a_6_n14# addersubtractor_0/fulladder_2/XOR_1/NAND_2/in1 0.12fF
C597 vdd comparator_0/XNOR_0/XOR_0/NAND_3/w_0_0# 0.05fF
C598 addersubtractor_0/fulladder_0/XOR_0/NAND_1/w_0_0# addersubtractor_0/fulladder_0/XOR_0/NAND_3/in1 0.03fF
C599 vdd enableblock_2/enable1_0/AND_3/not_0/w_0_0# 0.05fF
C600 AND_2/in1 comparator_0/NOR_0/w_32_0# 0.06fF
C601 comparator_0/XNOR_0/XOR_0/NAND_2/in1 comparator_0/XNOR_0/XOR_0/NAND_0/a_6_n14# 0.12fF
C602 comparator_0/XNOR_0/out comparator_0/threeinputAND_0/threeinputNAND_0/w_63_0# 0.06fF
C603 vdd addersubtractor_0/XOR_3/NAND_3/in1 0.25fF
C604 addersubtractor_0/XOR_0/out addersubtractor_0/XOR_0/NAND_3/a_6_n14# 0.12fF
C605 vdd comparator_0/XNOR_2/XOR_0/NAND_3/w_0_0# 0.05fF
C606 gnd comparator_0/XNOR_2/not_0/in 0.03fF
C607 twotofourdecoder_0/AND_3/NAND_0/w_0_0# twotofourdecoder_0/AND_3/not_0/in 0.03fF
C608 XOR_0/NAND_3/in1 XOR_0/NAND_1/a_6_n14# 0.12fF
C609 gnd comparator_0/XNOR_3/XOR_0/NAND_2/in1 0.15fF
C610 vdd comparator_0/not_3/out 0.07fF
C611 vdd and1 0.20fF
C612 comparator_0/fourinputOR_0/in2 comparator_0/XNOR_2/out 0.13fF
C613 addersubtractor_0/fulladder_0/XOR_1/NAND_2/a_6_n14# addersubtractor_0/fulladder_0/XOR_1/NAND_3/in2 0.12fF
C614 vdd comparator_0/fourinputAND_1/not_0/w_0_0# 0.05fF
C615 vdd comparator_0/XNOR_3/XOR_0/NAND_3/w_0_0# 0.05fF
C616 gnd comparator_0/XNOR_3/not_0/in 0.03fF
C617 XOR_0/NAND_2/w_0_0# XOR_0/NAND_3/in2 0.03fF
C618 vdd comparator_0/not_0/out 0.07fF
C619 gnd B1 0.86fF
C620 S0 B0 0.17fF
C621 enableblock_2/En enableblock_2/enable1_0/AND_1/NAND_0/w_0_0# 0.06fF
C622 andblock_0/AND_3/not_0/in andblock_0/AND_3/NAND_0/a_6_n14# 0.12fF
C623 comparator_0/fourinputAND_1/fourinputNAND_0/w_0_0# comparator_0/XNOR_3/out 0.06fF
C624 addersubtractor_0/fulladder_0/XOR_0/NAND_2/a_6_n14# addersubtractor_0/fulladder_0/XOR_0/NAND_3/in2 0.12fF
C625 enableblock_0/A_out3 gnd 1.67fF
C626 gnd twotofourdecoder_0/AND_3/not_0/in 0.04fF
C627 addersubtractor_0/XOR_2/NAND_2/in1 addersubtractor_0/XOR_2/NAND_2/w_0_0# 0.06fF
C628 addersubtractor_0/fulladder_1/XOR_0/NAND_2/in1 gnd 0.15fF
C629 vdd addersubtractor_0/fulladder_1/AND_0/NAND_0/w_0_0# 0.05fF
C630 comparator_0/fourinputAND_0/fourinputNAND_0/w_100_0# comparator_0/fourinputAND_0/not_0/in 0.03fF
C631 addersubtractor_0/fulladder_1/XOR_1/NAND_2/w_32_0# addersubtractor_0/fulladder_1/XOR_1/NAND_3/in2 0.03fF
C632 addersubtractor_0/fulladder_1/OR_0/in2 addersubtractor_0/fulladder_1/OR_0/NOR_0/w_32_0# 0.06fF
C633 enableblock_2/enable1_0/AND_2/NAND_0/w_32_0# enableblock_2/enable1_0/AND_2/not_0/in 0.03fF
C634 S0 enableblock_0/A_out0 0.06fF
C635 vdd addersubtractor_0/fulladder_2/AND_1/NAND_0/w_0_0# 0.05fF
C636 comparator_0/XNOR_0/out comparator_0/B1 0.06fF
C637 addersubtractor_0/fulladder_2/AND_0/not_0/in gnd 0.04fF
C638 addersubtractor_0/fulladder_0/OR_0/NOR_0/a_13_6# vdd 0.21fF
C639 addersubtractor_0/fulladder_0/OR_0/in1 gnd 0.30fF
C640 vdd enableblock_2/enable1_1/AND_1/not_0/in 0.29fF
C641 enableblock_2/enable1_0/AND_3/not_0/w_0_0# andblock_0/B2 0.03fF
C642 addersubtractor_0/fulladder_3/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_3/XOR_1/NAND_0/w_0_0# 0.03fF
C643 addersubtractor_0/XOR_0/out vdd 0.32fF
C644 comparator_0/XNOR_0/out comparator_0/B0 0.06fF
C645 comparator_0/fourinputAND_0/not_0/in comparator_0/fourinputAND_0/fourinputNAND_0/a_6_n14# 0.11fF
C646 addersubtractor_0/fulladder_1/XOR_0/NAND_2/w_32_0# addersubtractor_0/fulladder_1/XOR_0/NAND_3/in2 0.03fF
C647 vdd addersubtractor_0/fulladder_1/XOR_0/NAND_0/w_32_0# 0.05fF
C648 addersubtractor_0/XOR_1/NAND_2/w_32_0# addersubtractor_0/XOR_1/NAND_3/in2 0.03fF
C649 comparator_0/XNOR_1/XOR_0/NAND_0/w_32_0# comparator_0/B2 0.06fF
C650 vdd comparator_0/XNOR_1/XOR_0/NAND_0/w_0_0# 0.05fF
C651 vdd addersubtractor_0/fulladder_1/XOR_1/NAND_0/w_32_0# 0.05fF
C652 addersubtractor_0/fulladder_1/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_1/XOR_1/NAND_0/w_32_0# 0.03fF
C653 comparator_0/AND_0/not_0/w_0_0# comparator_0/AND_0/out 0.03fF
C654 comparator_0/fiveinputAND_0/fiveinputNAND_0/w_133_0# comparator_0/XNOR_2/out 0.06fF
C655 addersubtractor_0/XOR_1/NAND_2/in1 addersubtractor_0/XOR_1/NAND_0/a_6_n14# 0.12fF
C656 addersubtractor_0/XOR_2/out gnd 0.56fF
C657 comparator_0/XNOR_0/out comparator_0/XNOR_0/not_0/w_0_0# 0.03fF
C658 A0 B3 0.19fF
C659 addersubtractor_0/XOR_3/NAND_3/in1 addersubtractor_0/XOR_3/NAND_1/w_0_0# 0.03fF
C660 vdd addersubtractor_0/fulladder_3/AND_0/NAND_0/w_32_0# 0.05fF
C661 enableblock_0/enable1_0/AND_2/not_0/w_0_0# enableblock_0/enable1_0/AND_2/not_0/in 0.06fF
C662 enableblock_1/enable1_0/AND_1/not_0/w_0_0# comparator_0/B3 0.03fF
C663 addersubtractor_0/fulladder_2/XOR_1/in2 addersubtractor_0/fulladder_2/XOR_1/NAND_2/w_32_0# 0.06fF
C664 vdd addersubtractor_0/fulladder_2/OR_0/NOT_0/w_0_0# 0.05fF
C665 comparator_0/threeinputAND_0/threeinputNAND_0/a_45_n14# comparator_0/A2 0.18fF
C666 comparator_0/XNOR_2/out comparator_0/B1 0.84fF
C667 comparator_0/XNOR_2/XOR_0/NAND_2/in1 comparator_0/XNOR_2/XOR_0/NAND_0/a_6_n14# 0.12fF
C668 comparator_0/fourinputOR_0/fourinputNOR_0/w_32_0# comparator_0/fourinputOR_0/in2 0.06fF
C669 B1 enableblock_2/enable1_1/AND_1/NAND_0/w_32_0# 0.06fF
C670 gnd AND_0/in1 0.08fF
C671 vdd addersubtractor_0/fulladder_3/AND_1/not_0/in 0.29fF
C672 comparator_0/XNOR_1/not_0/w_0_0# comparator_0/XNOR_1/not_0/in 0.06fF
C673 enableblock_0/enable1_1/AND_0/NAND_0/w_0_0# A2 0.06fF
C674 addersubtractor_0/fulladder_3/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_3/XOR_1/NAND_1/a_6_n14# 0.12fF
C675 AND_2/in2 twotofourdecoder_0/AND_1/not_0/in 0.02fF
C676 comparator_0/XNOR_2/out comparator_0/B0 0.06fF
C677 comparator_0/fiveinputAND_0/fiveinputNAND_0/a_45_n14# comparator_0/fiveinputAND_0/fiveinputNAND_0/a_76_n14# 0.04fF
C678 enableblock_1/enable1_1/AND_2/NAND_0/w_32_0# enableblock_1/enable1_1/AND_2/not_0/in 0.03fF
C679 andblock_0/AND_1/not_0/w_0_0# andblock_0/AND_1/not_0/in 0.06fF
C680 twotofourdecoder_0/AND_2/NAND_0/w_32_0# twotofourdecoder_0/not_1/out 0.06fF
C681 vdd addersubtractor_0/fulladder_3/OR_0/NOR_0/w_0_0# 0.05fF
C682 vdd enableblock_1/enable1_1/AND_3/NAND_0/w_0_0# 0.05fF
C683 addersubtractor_0/fulladder_2/OR_0/NOR_0/a_13_6# addersubtractor_0/fulladder_2/OR_0/NOR_0/w_32_0# 0.03fF
C684 addersubtractor_0/fulladder_1/AND_0/not_0/in addersubtractor_0/fulladder_1/OR_0/in2 0.02fF
C685 andblock_0/AND_1/NAND_0/w_0_0# andblock_0/AND_1/not_0/in 0.03fF
C686 vdd comparator_0/XNOR_0/XOR_0/NAND_0/w_32_0# 0.05fF
C687 addersubtractor_0/fulladder_3/XOR_0/NAND_3/in1 addersubtractor_0/fulladder_3/XOR_0/NAND_1/a_6_n14# 0.12fF
C688 comparator_0/B2 comparator_0/XNOR_1/XOR_0/NAND_2/w_32_0# 0.06fF
C689 vdd enableblock_2/enable1_0/AND_2/NAND_0/w_32_0# 0.05fF
C690 vdd addersubtractor_0/XOR_3/NAND_2/in1 0.25fF
C691 addersubtractor_0/fulladder_3/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_3/XOR_1/NAND_2/w_0_0# 0.06fF
C692 twotofourdecoder_0/not_0/out twotofourdecoder_0/not_0/w_0_0# 0.03fF
C693 addersubtractor_0/fulladder_3/XOR_1/in2 addersubtractor_0/fulladder_3/XOR_1/NAND_0/w_32_0# 0.06fF
C694 vdd comparator_0/XNOR_2/XOR_0/NAND_0/w_32_0# 0.05fF
C695 comparator_0/XNOR_0/XOR_0/NAND_2/in1 comparator_0/XNOR_0/XOR_0/NAND_2/w_0_0# 0.06fF
C696 comparator_0/XNOR_1/XOR_0/NAND_3/in1 comparator_0/XNOR_1/XOR_0/NAND_1/a_6_n14# 0.12fF
C697 twotofourdecoder_0/AND_1/NAND_0/a_6_n14# twotofourdecoder_0/AND_1/not_0/in 0.12fF
C698 vdd enableblock_2/enable1_1/AND_0/NAND_0/w_0_0# 0.05fF
C699 vdd comparator_0/XNOR_3/XOR_0/NAND_0/w_32_0# 0.05fF
C700 vdd enableblock_0/enable1_0/AND_1/NAND_0/w_0_0# 0.05fF
C701 gnd AND_2/NAND_0/a_6_n14# 0.57fF
C702 addersubtractor_0/fulladder_0/OR_0/NOR_0/a_13_6# addersubtractor_0/fulladder_0/OR_0/NOR_0/w_0_0# 0.03fF
C703 AND_0/NAND_0/w_32_0# OR_0/out 0.06fF
C704 vdd lesser 0.43fF
C705 addersubtractor_0/fulladder_1/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_1/XOR_0/NAND_0/w_0_0# 0.03fF
C706 addersubtractor_0/fulladder_0/XOR_1/NAND_3/in1 gnd 0.11fF
C707 vdd addersubtractor_0/fulladder_0/XOR_1/NAND_1/w_0_0# 0.05fF
C708 comparator_0/XNOR_0/XOR_0/NAND_3/in1 comparator_0/XNOR_0/XOR_0/NAND_1/a_6_n14# 0.12fF
C709 A2 B3 4.40fF
C710 gnd enableblock_1/enable1_0/AND_3/NAND_0/a_6_n14# 0.57fF
C711 vdd enableblock_1/enable1_0/AND_2/not_0/w_0_0# 0.05fF
C712 addersubtractor_0/fulladder_0/XOR_0/NAND_3/in1 gnd 0.11fF
C713 addersubtractor_0/fulladder_0/XOR_0/NAND_1/w_0_0# vdd 0.05fF
C714 enableblock_0/enable1_0/AND_1/NAND_0/a_6_n14# enableblock_0/enable1_0/AND_1/not_0/in 0.12fF
C715 comparator_0/A3 comparator_0/B3 0.38fF
C716 A0 enableblock_2/enable1_1/AND_2/NAND_0/w_0_0# 0.06fF
C717 enableblock_0/A_out1 addersubtractor_0/XOR_1/out 0.11fF
C718 addersubtractor_0/fulladder_1/XOR_1/NAND_1/a_6_n14# gnd 0.57fF
C719 vdd XOR_0/NAND_1/w_32_0# 0.05fF
C720 addersubtractor_0/fulladder_2/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_2/XOR_0/NAND_0/w_32_0# 0.03fF
C721 addersubtractor_0/fulladder_2/AND_1/not_0/w_0_0# addersubtractor_0/fulladder_2/AND_1/not_0/in 0.06fF
C722 vdd addersubtractor_0/fulladder_1/XOR_1/NAND_1/w_32_0# 0.05fF
C723 addersubtractor_0/fulladder_1/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_1/XOR_1/NAND_1/w_32_0# 0.06fF
C724 enableblock_2/enable1_1/AND_3/NAND_0/w_0_0# enableblock_2/enable1_1/AND_3/not_0/in 0.03fF
C725 vdd andblock_0/A0 0.20fF
C726 enableblock_0/enable1_0/AND_1/not_0/w_0_0# enableblock_0/A_out2 0.03fF
C727 addersubtractor_0/fulladder_1/XOR_0/NAND_1/a_6_n14# gnd 0.57fF
C728 comparator_0/XNOR_2/XOR_0/NAND_3/in1 comparator_0/XNOR_2/XOR_0/NAND_1/a_6_n14# 0.12fF
C729 addersubtractor_0/XOR_2/NAND_3/in1 addersubtractor_0/XOR_2/NAND_3/w_0_0# 0.06fF
C730 vdd addersubtractor_0/fulladder_1/XOR_0/NAND_1/w_32_0# 0.05fF
C731 gnd enableblock_0/enable1_1/AND_1/not_0/in 0.04fF
C732 A0 enableblock_0/enable1_0/AND_0/NAND_0/w_0_0# 0.06fF
C733 comparator_0/A1 comparator_0/B1 0.95fF
C734 addersubtractor_0/XOR_2/NAND_0/w_0_0# addersubtractor_0/XOR_2/NAND_2/in1 0.03fF
C735 enableblock_0/enable1_1/AND_2/NAND_0/a_6_n14# enableblock_0/enable1_1/AND_2/not_0/in 0.12fF
C736 gnd and0 0.08fF
C737 comparator_0/AND_0/out comparator_0/fourinputOR_0/in2 1.17fF
C738 enableblock_0/enable1_1/AND_0/NAND_0/a_6_n14# enableblock_0/enable1_1/AND_0/not_0/in 0.12fF
C739 A3 B3 0.23fF
C740 OR_0/in2 OR_0/NOT_0/in 0.26fF
C741 comparator_0/XNOR_3/XOR_0/NAND_3/in1 comparator_0/XNOR_3/XOR_0/NAND_1/a_6_n14# 0.12fF
C742 enableblock_1/enable1_0/AND_0/not_0/w_0_0# enableblock_1/enable1_0/AND_0/not_0/in 0.06fF
C743 addersubtractor_0/XOR_0/NAND_2/in1 addersubtractor_0/XOR_0/NAND_0/w_0_0# 0.03fF
C744 vdd comparator_0/AND_0/not_0/in 0.29fF
C745 OR_0/out enableblock_0/enable1_0/AND_3/NAND_0/w_0_0# 0.06fF
C746 A1 enableblock_0/enable1_0/AND_2/NAND_0/w_0_0# 0.06fF
C747 comparator_0/A0 comparator_0/B0 0.13fF
C748 comparator_0/not_1/w_0_0# comparator_0/B2 0.06fF
C749 vdd andblock_0/AND_0/not_0/in 0.29fF
C750 comparator_0/XNOR_2/XOR_0/NAND_2/in1 comparator_0/XNOR_2/XOR_0/NAND_2/w_0_0# 0.06fF
C751 enableblock_1/enable1_0/AND_0/NAND_0/a_6_n14# A3 0.07fF
C752 gnd enableblock_0/enable1_0/AND_1/NAND_0/a_6_n14# 0.57fF
C753 vdd addersubtractor_0/fulladder_2/C 0.18fF
C754 vdd enableblock_2/enable1_1/AND_0/not_0/in 0.29fF
C755 vdd enableblock_0/enable1_0/AND_0/not_0/w_0_0# 0.05fF
C756 enableblock_0/enable1_0/AND_3/NAND_0/w_32_0# enableblock_0/enable1_0/AND_3/not_0/in 0.03fF
C757 gnd addersubtractor_0/XOR_3/NAND_3/a_6_n14# 0.57fF
C758 vdd addersubtractor_0/XOR_3/NAND_3/w_32_0# 0.05fF
C759 addersubtractor_0/fulladder_3/AND_1/not_0/w_0_0# addersubtractor_0/fulladder_3/OR_0/in1 0.03fF
C760 AND_2/in2 OR_0/in2 1.07fF
C761 comparator_0/A2 comparator_0/XNOR_1/XOR_0/NAND_1/w_0_0# 0.06fF
C762 comparator_0/XNOR_3/out comparator_0/XNOR_3/not_0/w_0_0# 0.03fF
C763 OR_0/in2 twotofourdecoder_0/AND_2/not_0/in 0.02fF
C764 vdd enableblock_1/enable1_1/AND_3/not_0/in 0.29fF
C765 gnd enableblock_2/enable1_0/AND_2/not_0/in 0.04fF
C766 addersubtractor_0/XOR_1/out addersubtractor_0/XOR_1/NAND_3/w_32_0# 0.03fF
C767 and0 andblock_0/AND_3/not_0/w_0_0# 0.03fF
C768 twotofourdecoder_0/AND_0/NAND_0/w_32_0# S1 0.06fF
C769 gnd addersubtractor_0/XOR_2/NAND_1/a_6_n14# 0.57fF
C770 vdd addersubtractor_0/XOR_2/NAND_1/w_32_0# 0.05fF
C771 comparator_0/A3 comparator_0/XNOR_0/XOR_0/NAND_0/w_0_0# 0.06fF
C772 vdd enableblock_2/enable1_1/AND_0/not_0/w_0_0# 0.05fF
C773 enableblock_1/enable1_0/AND_3/not_0/w_0_0# enableblock_1/enable1_0/AND_3/not_0/in 0.06fF
C774 vdd andblock_0/AND_2/not_0/w_0_0# 0.05fF
C775 vdd enableblock_0/enable1_0/AND_1/not_0/in 0.29fF
C776 andblock_0/A2 andblock_0/AND_1/NAND_0/a_6_n14# 0.02fF
C777 vdd enableblock_1/enable1_0/AND_1/NAND_0/w_32_0# 0.05fF
C778 gnd addersubtractor_0/XOR_0/NAND_3/a_6_n14# 0.57fF
C779 XOR_0/NAND_0/a_6_n14# XOR_0/NAND_2/in1 0.12fF
C780 comparator_0/XNOR_0/out comparator_0/XNOR_1/out 1.10fF
C781 enableblock_1/enable1_1/AND_3/NAND_0/w_32_0# B0 0.06fF
C782 enableblock_1/enable1_0/AND_3/NAND_0/w_32_0# B2 0.06fF
C783 enableblock_1/enable1_0/AND_1/NAND_0/w_32_0# B3 0.06fF
C784 vdd addersubtractor_0/XOR_0/NAND_3/w_32_0# 0.05fF
C785 enableblock_0/A_out1 addersubtractor_0/fulladder_1/XOR_0/NAND_1/w_0_0# 0.06fF
C786 comparator_0/not_0/out comparator_0/not_0/w_0_0# 0.03fF
C787 comparator_0/A1 comparator_0/XNOR_2/XOR_0/NAND_0/w_0_0# 0.06fF
C788 gnd andblock_0/A3 0.10fF
C789 AND_2/in2 enableblock_1/enable1_1/AND_2/NAND_0/w_32_0# 0.06fF
C790 AND_2/NAND_0/w_0_0# AND_2/not_0/in 0.03fF
C791 addersubtractor_0/fulladder_1/XOR_1/NAND_3/w_32_0# addersubtractor_0/fulladder_1/XOR_1/NAND_3/in2 0.06fF
C792 vdd twotofourdecoder_0/AND_3/NAND_0/w_0_0# 0.05fF
C793 vdd addersubtractor_0/XOR_2/NAND_0/w_32_0# 0.05fF
C794 enableblock_1/enable1_1/AND_1/NAND_0/a_6_n14# enableblock_1/enable1_1/AND_1/not_0/in 0.12fF
C795 gnd enableblock_1/enable1_1/AND_0/NAND_0/a_6_n14# 0.57fF
C796 addersubtractor_0/fulladder_2/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_2/XOR_0/NAND_1/w_32_0# 0.06fF
C797 gnd twotofourdecoder_0/AND_0/NAND_0/a_6_n14# 0.57fF
C798 A1 enableblock_2/En 0.13fF
C799 enableblock_1/enable1_0/AND_3/not_0/w_0_0# comparator_0/B2 0.03fF
C800 addersubtractor_0/fulladder_0/XOR_1/NAND_0/a_6_n14# gnd 0.57fF
C801 addersubtractor_0/fulladder_0/AND_0/not_0/w_0_0# addersubtractor_0/fulladder_0/OR_0/in2 0.03fF
C802 vdd enableblock_2/enable1_1/AND_3/not_0/w_0_0# 0.05fF
C803 vdd enableblock_2/enable1_0/AND_0/NAND_0/w_0_0# 0.05fF
C804 enableblock_0/enable1_1/AND_1/NAND_0/w_0_0# enableblock_0/enable1_1/AND_1/not_0/in 0.03fF
C805 comparator_0/A0 comparator_0/XNOR_3/XOR_0/NAND_0/w_0_0# 0.06fF
C806 addersubtractor_0/fulladder_1/XOR_0/NAND_3/w_32_0# addersubtractor_0/fulladder_1/XOR_0/NAND_3/in2 0.06fF
C807 comparator_0/fiveinputAND_0/fiveinputNAND_0/w_63_0# comparator_0/XNOR_1/out 0.06fF
C808 enableblock_2/enable1_0/AND_3/NAND_0/a_6_n14# enableblock_2/enable1_0/AND_3/not_0/in 0.12fF
C809 adder1 addersubtractor_0/fulladder_1/XOR_1/NAND_3/a_6_n14# 0.12fF
C810 gnd andblock_0/AND_3/not_0/in 0.04fF
C811 addersubtractor_0/XOR_1/NAND_3/w_32_0# addersubtractor_0/XOR_1/NAND_3/in2 0.06fF
C812 vdd addersubtractor_0/fulladder_1/XOR_1/NAND_3/in2 0.25fF
C813 comparator_0/fourinputAND_0/fourinputNAND_0/a_76_n14# comparator_0/XNOR_1/out 0.23fF
C814 vdd enableblock_1/enable1_1/AND_0/NAND_0/w_32_0# 0.05fF
C815 addersubtractor_0/fulladder_3/OR_0/in2 addersubtractor_0/fulladder_3/OR_0/NOT_0/in 0.26fF
C816 vdd gnd 7.13fF
C817 andblock_0/AND_3/not_0/in andblock_0/AND_3/NAND_0/w_32_0# 0.03fF
C818 comparator_0/fourinputAND_1/fourinputNAND_0/w_100_0# comparator_0/fourinputAND_1/not_0/in 0.03fF
C819 addersubtractor_0/fulladder_1/XOR_1/NAND_2/in1 gnd 0.15fF
C820 vdd addersubtractor_0/fulladder_1/XOR_0/NAND_3/in2 0.25fF
C821 comparator_0/XNOR_2/out comparator_0/XNOR_1/out 0.21fF
C822 gnd B3 0.91fF
C823 addersubtractor_0/fulladder_1/XOR_1/in2 addersubtractor_0/fulladder_1/XOR_0/NAND_3/a_6_n14# 0.12fF
C824 comparator_0/fourinputOR_0/fourinputNOR_0/w_0_0# comparator_0/AND_0/out 0.06fF
C825 enableblock_2/En enableblock_2/enable1_1/AND_1/NAND_0/w_0_0# 0.06fF
C826 vdd addersubtractor_0/fulladder_3/AND_0/not_0/w_0_0# 0.05fF
C827 addersubtractor_0/fulladder_0/AND_0/not_0/in vdd 0.29fF
C828 S0 B2 0.20fF
C829 vdd andblock_0/AND_3/NAND_0/w_32_0# 0.05fF
C830 gnd comparator_0/fourinputAND_1/fourinputNAND_0/a_76_n14# 0.04fF
C831 twotofourdecoder_0/AND_1/not_0/w_0_0# twotofourdecoder_0/AND_1/not_0/in 0.06fF
C832 vdd AND_2/not_0/w_0_0# 0.05fF
C833 addersubtractor_0/fulladder_2/XOR_1/NAND_3/w_32_0# adder2 0.03fF
C834 gnd enableblock_1/enable1_0/AND_0/NAND_0/a_6_n14# 0.57fF
C835 gnd comparator_0/XNOR_1/XOR_0/NAND_0/a_6_n14# 0.57fF
C836 twotofourdecoder_0/AND_0/not_0/in twotofourdecoder_0/AND_0/NAND_0/w_0_0# 0.03fF
C837 vdd addersubtractor_0/fulladder_0/XOR_1/NAND_0/w_0_0# 0.05fF
C838 enableblock_2/En S1 0.07fF
C839 comparator_0/fourinputAND_1/not_0/in comparator_0/fourinputAND_1/fourinputNAND_0/a_6_n14# 0.11fF
C840 comparator_0/not_3/w_0_0# comparator_0/not_3/out 0.03fF
C841 vdd and3 0.20fF
C842 S0 enableblock_0/B_out0 0.06fF
C843 gnd comparator_0/threeinputAND_0/threeinputNAND_0/a_6_n14# 0.47fF
C844 addersubtractor_0/fulladder_2/XOR_0/NAND_3/w_32_0# addersubtractor_0/fulladder_2/XOR_1/in2 0.03fF
C845 enableblock_1/enable1_0/AND_1/NAND_0/w_32_0# enableblock_1/enable1_0/AND_1/not_0/in 0.03fF
C846 comparator_0/fiveinputAND_0/not_0/w_0_0# comparator_0/fiveinputAND_0/not_0/in 0.06fF
C847 gnd enableblock_0/enable1_1/AND_0/not_0/in 0.04fF
C848 vdd addersubtractor_0/XOR_0/NAND_1/w_32_0# 0.05fF
C849 gnd comparator_0/XNOR_1/XOR_0/NAND_3/in2 0.07fF
C850 gnd comparator_0/not_2/out 0.08fF
C851 vdd adder3 0.25fF
C852 S0 addersubtractor_0/XOR_0/NAND_0/w_32_0# 0.06fF
C853 vdd addersubtractor_0/fulladder_2/OR_0/NOR_0/w_32_0# 0.03fF
C854 enableblock_0/enable1_0/AND_0/NAND_0/w_32_0# OR_0/out 0.06fF
C855 enableblock_1/enable1_1/AND_0/NAND_0/w_0_0# A1 0.06fF
C856 addersubtractor_0/XOR_3/out addersubtractor_0/XOR_3/NAND_3/w_0_0# 0.03fF
C857 vdd addersubtractor_0/fulladder_3/XOR_1/in2 0.47fF
C858 andblock_0/AND_3/not_0/w_0_0# andblock_0/AND_3/not_0/in 0.06fF
C859 gnd comparator_0/XNOR_0/XOR_0/NAND_3/in2 0.07fF
C860 gnd andblock_0/B2 0.38fF
C861 vdd andblock_0/AND_3/not_0/w_0_0# 0.05fF
C862 vdd comparator_0/XNOR_1/not_0/in 0.25fF
C863 comparator_0/threeinputAND_0/threeinputNAND_0/w_0_0# comparator_0/not_1/out 0.06fF
C864 S1 twotofourdecoder_0/AND_1/NAND_0/w_0_0# 0.06fF
C865 enableblock_2/enable1_0/AND_1/NAND_0/w_32_0# enableblock_2/enable1_0/AND_1/not_0/in 0.03fF
C866 enableblock_1/enable1_1/AND_3/NAND_0/a_6_n14# enableblock_1/enable1_1/AND_3/not_0/in 0.12fF
C867 gnd comparator_0/XNOR_2/XOR_0/NAND_3/in2 0.07fF
C868 gnd XOR_0/in1 0.88fF
C869 vdd comparator_0/fiveinputAND_0/fiveinputNAND_0/w_100_0# 0.05fF
C870 gnd addersubtractor_0/XOR_0/NAND_2/a_6_n14# 0.59fF
C871 vdd comparator_0/XNOR_0/not_0/in 0.25fF
C872 vdd comparator_0/fourinputOR_0/in4 0.93fF
C873 addersubtractor_0/fulladder_1/AND_0/NAND_0/a_6_n14# gnd 0.57fF
C874 AND_2/in2 greater 0.06fF
C875 S1 twotofourdecoder_0/not_1/w_0_0# 0.06fF
C876 vdd enableblock_2/enable1_1/AND_1/NAND_0/w_32_0# 0.05fF
C877 gnd comparator_0/XNOR_3/XOR_0/NAND_3/in2 0.07fF
C878 addersubtractor_0/fulladder_1/XOR_1/NAND_1/w_0_0# addersubtractor_0/fulladder_1/XOR_1/NAND_3/in1 0.03fF
C879 AND_2/in2 B2 0.06fF
C880 vdd comparator_0/XNOR_2/not_0/in 0.25fF
C881 enableblock_1/enable1_1/AND_1/not_0/w_0_0# comparator_0/B1 0.03fF
C882 S0 OR_0/out 1.74fF
C883 vdd comparator_0/XNOR_3/XOR_0/NAND_2/in1 0.25fF
C884 gnd comparator_0/fiveinputAND_0/fiveinputNAND_0/a_113_n14# 0.04fF
C885 gnd enableblock_1/enable1_0/AND_1/not_0/in 0.04fF
C886 comparator_0/AND_0/NAND_0/w_32_0# comparator_0/AND_0/not_0/in 0.03fF
C887 addersubtractor_0/fulladder_0/AND_1/not_0/in gnd 0.04fF
C888 andblock_0/A0 enableblock_2/enable1_1/AND_2/not_0/in 0.02fF
C889 AND_2/NAND_0/w_32_0# AND_2/not_0/in 0.03fF
C890 addersubtractor_0/fulladder_3/XOR_1/NAND_0/a_6_n14# addersubtractor_0/fulladder_3/XOR_1/NAND_2/in1 0.12fF
C891 comparator_0/fourinputAND_0/fourinputNAND_0/w_32_0# comparator_0/fourinputAND_0/not_0/in 0.03fF
C892 addersubtractor_0/fulladder_2/OR_0/in2 gnd 0.36fF
C893 addersubtractor_0/fulladder_1/XOR_0/NAND_1/w_0_0# addersubtractor_0/fulladder_1/XOR_0/NAND_3/in1 0.03fF
C894 comparator_0/XNOR_0/out comparator_0/XNOR_2/out 0.51fF
C895 vdd comparator_0/XNOR_3/not_0/in 0.25fF
C896 vdd comparator_0/fourinputOR_0/fourinputNOR_0/w_64_0# 0.03fF
C897 enableblock_1/enable1_0/AND_0/NAND_0/w_32_0# AND_2/in2 0.06fF
C898 vdd addersubtractor_0/fulladder_0/XOR_1/NAND_2/w_0_0# 0.05fF
C899 comparator_0/fourinputAND_1/fourinputNAND_0/w_0_0# comparator_0/fourinputAND_1/not_0/in 0.03fF
C900 B1 B3 0.19fF
C901 addersubtractor_0/fulladder_0/XOR_0/NAND_2/w_0_0# vdd 0.05fF
C902 XOR_0/NAND_1/w_32_0# XOR_0/NAND_2/in1 0.06fF
C903 comparator_0/fiveinputAND_0/not_0/in comparator_0/fiveinputAND_0/fiveinputNAND_0/a_6_n14# 0.11fF
C904 gnd comparator_0/fourinputOR_0/not_0/in 0.94fF
C905 vdd enableblock_2/enable1_1/AND_2/NAND_0/w_32_0# 0.05fF
C906 enableblock_0/A_out3 vdd 0.43fF
C907 vdd addersubtractor_0/fulladder_1/XOR_0/NAND_2/in1 0.25fF
C908 vdd twotofourdecoder_0/AND_3/not_0/in 0.29fF
C909 addersubtractor_0/fulladder_1/XOR_1/NAND_2/a_6_n14# addersubtractor_0/fulladder_1/XOR_1/NAND_3/in2 0.12fF
C910 comparator_0/A1 comparator_0/XNOR_1/out 0.06fF
C911 enableblock_2/enable1_0/AND_2/NAND_0/w_0_0# enableblock_2/enable1_0/AND_2/not_0/in 0.03fF
C912 comparator_0/fourinputOR_0/fourinputNOR_0/a_77_6# comparator_0/fourinputOR_0/fourinputNOR_0/w_97_0# 0.03fF
C913 addersubtractor_0/fulladder_1/XOR_1/NAND_2/a_6_n14# gnd 0.59fF
C914 vdd addersubtractor_0/fulladder_1/XOR_1/NAND_2/w_32_0# 0.05fF
C915 vdd OR_0/NOT_0/w_0_0# 0.05fF
C916 vdd addersubtractor_0/fulladder_2/AND_0/not_0/in 0.29fF
C917 vdd comparator_0/XNOR_1/not_0/w_0_0# 0.05fF
C918 addersubtractor_0/fulladder_0/OR_0/in1 vdd 0.12fF
C919 addersubtractor_0/fulladder_1/XOR_0/NAND_2/a_6_n14# gnd 0.59fF
C920 vdd addersubtractor_0/fulladder_1/XOR_0/NAND_2/w_32_0# 0.05fF
C921 OR_0/out OR_0/NOT_0/in 0.02fF
C922 comparator_0/A0 comparator_0/XNOR_1/out 0.10fF
C923 enableblock_0/B_out3 gnd 1.68fF
C924 addersubtractor_0/fulladder_1/XOR_0/NAND_2/a_6_n14# addersubtractor_0/fulladder_1/XOR_0/NAND_3/in2 0.12fF
C925 vdd addersubtractor_0/fulladder_1/XOR_0/NAND_0/w_0_0# 0.05fF
C926 addersubtractor_0/fulladder_1/AND_1/NAND_0/a_6_n14# addersubtractor_0/fulladder_1/AND_1/not_0/in 0.12fF
C927 gnd addersubtractor_0/fulladder_3/XOR_0/NAND_2/in1 0.15fF
C928 addersubtractor_0/fulladder_1/AND_1/NAND_0/w_0_0# vdd 0.05fF
C929 vdd enableblock_0/enable1_1/AND_1/NAND_0/w_0_0# 0.05fF
C930 addersubtractor_0/XOR_2/NAND_1/w_32_0# addersubtractor_0/XOR_2/NAND_3/in1 0.03fF
C931 addersubtractor_0/XOR_1/NAND_2/a_6_n14# addersubtractor_0/XOR_1/NAND_3/in2 0.12fF
C932 vdd addersubtractor_0/fulladder_3/AND_0/NAND_0/w_0_0# 0.05fF
C933 addersubtractor_0/fulladder_2/XOR_1/NAND_2/w_32_0# addersubtractor_0/fulladder_2/XOR_1/NAND_3/in2 0.03fF
C934 addersubtractor_0/fulladder_2/OR_0/in2 addersubtractor_0/fulladder_2/OR_0/NOR_0/w_32_0# 0.06fF
C935 comparator_0/fiveinputAND_0/fiveinputNAND_0/w_0_0# comparator_0/not_3/out 0.06fF
C936 vdd addersubtractor_0/XOR_1/NAND_1/w_32_0# 0.05fF
C937 gnd addersubtractor_0/XOR_0/NAND_3/in1 0.11fF
C938 B0 A1 0.75fF
C939 addersubtractor_0/fulladder_2/OR_0/in1 gnd 0.30fF
C940 vdd addersubtractor_0/fulladder_2/OR_0/NOR_0/a_13_6# 0.21fF
C941 gnd enableblock_1/enable1_1/AND_3/NAND_0/a_6_n14# 0.57fF
C942 vdd addersubtractor_0/fulladder_3/XOR_0/NAND_0/w_32_0# 0.05fF
C943 vdd addersubtractor_0/XOR_2/out 0.32fF
C944 addersubtractor_0/fulladder_2/XOR_0/NAND_2/w_32_0# addersubtractor_0/fulladder_2/XOR_0/NAND_3/in2 0.03fF
C945 vdd enableblock_1/enable1_1/AND_2/not_0/w_0_0# 0.05fF
C946 addersubtractor_0/XOR_2/NAND_2/in1 addersubtractor_0/XOR_2/NAND_0/a_6_n14# 0.12fF
C947 enableblock_0/B_out1 enableblock_0/enable1_1/AND_2/not_0/in 0.02fF
C948 vdd addersubtractor_0/fulladder_3/XOR_1/NAND_0/w_32_0# 0.05fF
C949 addersubtractor_0/fulladder_2/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_2/XOR_1/NAND_0/w_32_0# 0.03fF
C950 comparator_0/fiveinputAND_0/fiveinputNAND_0/a_6_n14# comparator_0/fiveinputAND_0/fiveinputNAND_0/a_45_n14# 0.04fF
C951 twotofourdecoder_0/AND_2/NAND_0/w_32_0# twotofourdecoder_0/AND_2/not_0/in 0.03fF
C952 A0 enableblock_2/En 0.13fF
C953 vdd AND_0/in1 0.10fF
C954 comparator_0/fourinputOR_0/in4 comparator_0/fourinputOR_0/not_0/in 0.10fF
C955 addersubtractor_0/XOR_0/NAND_1/w_32_0# addersubtractor_0/XOR_0/NAND_3/in1 0.03fF
C956 addersubtractor_0/fulladder_0/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_0/XOR_0/NAND_0/a_6_n14# 0.12fF
C957 vdd comparator_0/XNOR_0/XOR_0/NAND_1/w_0_0# 0.05fF
C958 comparator_0/XNOR_3/XOR_0/NAND_2/in1 comparator_0/XNOR_3/XOR_0/NAND_1/w_32_0# 0.06fF
C959 comparator_0/fourinputOR_0/fourinputNOR_0/w_64_0# comparator_0/fourinputOR_0/fourinputNOR_0/a_45_6# 0.03fF
C960 enableblock_1/enable1_1/AND_2/NAND_0/w_0_0# enableblock_1/enable1_1/AND_2/not_0/in 0.03fF
C961 addersubtractor_0/fulladder_3/XOR_1/in2 addersubtractor_0/fulladder_3/XOR_1/NAND_2/w_32_0# 0.06fF
C962 B0 S1 0.06fF
C963 comparator_0/XNOR_0/out comparator_0/A3 0.01fF
C964 vdd comparator_0/XNOR_2/XOR_0/NAND_1/w_0_0# 0.05fF
C965 addersubtractor_0/fulladder_0/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_0/XOR_1/NAND_3/w_0_0# 0.06fF
C966 enableblock_2/enable1_1/AND_1/not_0/w_0_0# enableblock_2/enable1_1/AND_1/not_0/in 0.06fF
C967 addersubtractor_0/fulladder_1/AND_0/not_0/in addersubtractor_0/fulladder_1/AND_0/NAND_0/w_32_0# 0.03fF
C968 addersubtractor_0/fulladder_0/XOR_0/NAND_0/w_32_0# addersubtractor_0/XOR_0/out 0.06fF
C969 comparator_0/XNOR_0/XOR_0/NAND_2/in1 comparator_0/XNOR_0/XOR_0/NAND_0/w_32_0# 0.03fF
C970 vdd enableblock_2/enable1_0/AND_2/NAND_0/w_0_0# 0.05fF
C971 comparator_0/XNOR_0/out comparator_0/A1 0.06fF
C972 vdd comparator_0/XNOR_3/XOR_0/NAND_1/w_0_0# 0.05fF
C973 gnd addersubtractor_0/XOR_2/NAND_3/in1 0.11fF
C974 addersubtractor_0/XOR_1/NAND_1/w_0_0# enableblock_0/A_out0 0.06fF
C975 S0 addersubtractor_0/XOR_1/NAND_2/w_32_0# 0.06fF
C976 addersubtractor_0/fulladder_0/XOR_0/NAND_3/in1 addersubtractor_0/fulladder_0/XOR_0/NAND_3/w_0_0# 0.06fF
C977 OR_0/out enableblock_0/enable1_1/AND_3/NAND_0/w_0_0# 0.06fF
C978 addersubtractor_0/fulladder_3/OR_0/NOR_0/a_13_6# addersubtractor_0/fulladder_3/OR_0/NOR_0/w_32_0# 0.03fF
C979 addersubtractor_0/fulladder_2/AND_0/not_0/in addersubtractor_0/fulladder_2/OR_0/in2 0.02fF
C980 addersubtractor_0/fulladder_0/AND_1/not_0/in addersubtractor_0/fulladder_0/OR_0/in1 0.02fF
C981 comparator_0/XNOR_0/out comparator_0/A0 0.06fF
C982 addersubtractor_0/XOR_1/NAND_2/in1 addersubtractor_0/XOR_1/NAND_0/w_0_0# 0.03fF
C983 vdd enableblock_0/enable1_0/AND_3/not_0/w_0_0# 0.05fF
C984 enableblock_2/En enableblock_2/enable1_0/AND_2/NAND_0/w_32_0# 0.06fF
C985 vdd addersubtractor_0/XOR_0/out 0.06fF
C986 gnd AND_0/not_0/in 0.04fF
C987 addersubtractor_0/fulladder_2/AND_1/NAND_0/w_0_0# addersubtractor_0/fulladder_2/AND_1/not_0/in 0.03fF
C988 addersubtractor_0/fulladder_0/OR_0/NOR_0/w_0_0# addersubtractor_0/fulladder_0/OR_0/in1 0.06fF
C989 addersubtractor_0/XOR_0/NAND_2/w_0_0# addersubtractor_0/XOR_0/NAND_3/in2 0.03fF
C990 OR_0/NOR_0/a_13_6# OR_0/NOR_0/w_0_0# 0.03fF
C991 vdd comparator_0/fourinputOR_0/not_0/w_0_0# 0.05fF
C992 vdd addersubtractor_0/fulladder_0/XOR_1/NAND_3/in1 0.25fF
C993 gnd OR_0/in1 0.11fF
C994 XOR_0/NAND_3/in1 XOR_0/NAND_1/w_32_0# 0.03fF
C995 gnd enableblock_2/enable1_1/AND_2/not_0/in 0.04fF
C996 addersubtractor_0/fulladder_0/XOR_0/NAND_3/in1 vdd 0.25fF
C997 addersubtractor_0/fulladder_1/OR_0/NOT_0/in gnd 0.60fF
C998 addersubtractor_0/fulladder_1/OR_0/NOR_0/a_13_6# addersubtractor_0/fulladder_1/OR_0/NOR_0/w_0_0# 0.03fF
C999 comparator_0/XNOR_2/out comparator_0/A1 0.11fF
C1000 S0 twotofourdecoder_0/not_1/out 0.13fF
C1001 addersubtractor_0/XOR_2/NAND_1/w_32_0# addersubtractor_0/XOR_2/NAND_2/in1 0.06fF
C1002 A2 enableblock_2/En 0.13fF
C1003 gnd addersubtractor_0/fulladder_2/XOR_1/NAND_3/in1 0.11fF
C1004 addersubtractor_0/fulladder_2/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_2/XOR_0/NAND_0/w_0_0# 0.03fF
C1005 vdd addersubtractor_0/fulladder_2/XOR_1/NAND_1/w_0_0# 0.05fF
C1006 gnd XOR_0/NAND_2/in1 0.15fF
C1007 comparator_0/XNOR_2/out comparator_0/A0 0.06fF
C1008 addersubtractor_0/fulladder_2/XOR_0/NAND_3/in1 gnd 0.11fF
C1009 addersubtractor_0/fulladder_1/AND_1/NAND_0/a_6_n14# addersubtractor_0/fulladder_0/C 0.07fF
C1010 vdd enableblock_0/enable1_1/AND_1/not_0/in 0.29fF
C1011 vdd addersubtractor_0/fulladder_2/XOR_0/NAND_1/w_0_0# 0.05fF
C1012 comparator_0/fourinputOR_0/fourinputNOR_0/a_13_6# comparator_0/fourinputOR_0/fourinputNOR_0/w_0_0# 0.03fF
C1013 and0 andblock_0/AND_3/not_0/in 0.02fF
C1014 enableblock_0/B_out3 addersubtractor_0/XOR_2/out 0.11fF
C1015 gnd addersubtractor_0/fulladder_3/XOR_1/NAND_1/a_6_n14# 0.57fF
C1016 vdd addersubtractor_0/fulladder_3/XOR_1/NAND_1/w_32_0# 0.05fF
C1017 vdd and0 0.10fF
C1018 addersubtractor_0/fulladder_3/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_3/XOR_0/NAND_0/w_32_0# 0.03fF
C1019 addersubtractor_0/fulladder_3/AND_1/not_0/w_0_0# addersubtractor_0/fulladder_3/AND_1/not_0/in 0.06fF
C1020 addersubtractor_0/fulladder_2/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_2/XOR_1/NAND_1/w_32_0# 0.06fF
C1021 gnd addersubtractor_0/fulladder_3/XOR_0/NAND_1/a_6_n14# 0.57fF
C1022 vdd addersubtractor_0/fulladder_3/XOR_0/NAND_1/w_32_0# 0.05fF
C1023 addersubtractor_0/fulladder_0/AND_1/NAND_0/a_6_n14# S0 0.07fF
C1024 comparator_0/AND_0/out comparator_0/XNOR_0/out 0.06fF
C1025 comparator_0/XNOR_2/XOR_0/NAND_2/in1 comparator_0/XNOR_2/XOR_0/NAND_0/w_32_0# 0.03fF
C1026 enableblock_0/B_out0 enableblock_0/enable1_1/AND_3/not_0/in 0.02fF
C1027 gnd comparator_0/XNOR_1/XOR_0/NAND_1/a_6_n14# 0.57fF
C1028 addersubtractor_0/XOR_2/NAND_0/w_32_0# addersubtractor_0/XOR_2/NAND_2/in1 0.03fF
C1029 vdd comparator_0/XNOR_1/XOR_0/NAND_1/w_32_0# 0.05fF
C1030 vdd andblock_0/AND_2/NAND_0/w_0_0# 0.05fF
C1031 A3 enableblock_2/En 0.13fF
C1032 gnd comparator_0/XNOR_0/XOR_0/NAND_1/a_6_n14# 0.57fF
C1033 addersubtractor_0/XOR_3/NAND_2/w_0_0# addersubtractor_0/XOR_3/NAND_3/in2 0.03fF
C1034 enableblock_0/enable1_0/AND_3/NAND_0/w_0_0# enableblock_0/enable1_0/AND_3/not_0/in 0.03fF
C1035 gnd comparator_0/XNOR_2/XOR_0/NAND_1/a_6_n14# 0.57fF
C1036 enableblock_1/enable1_0/AND_2/NAND_0/a_6_n14# enableblock_1/enable1_0/AND_2/not_0/in 0.12fF
C1037 gnd addersubtractor_0/XOR_2/NAND_2/in1 0.15fF
C1038 vdd addersubtractor_0/XOR_1/NAND_2/w_0_0# 0.05fF
C1039 A0 B0 0.15fF
C1040 addersubtractor_0/XOR_1/out addersubtractor_0/XOR_1/NAND_3/a_6_n14# 0.12fF
C1041 vdd enableblock_2/enable1_0/AND_2/not_0/in 0.29fF
C1042 gnd comparator_0/XNOR_3/XOR_0/NAND_1/a_6_n14# 0.57fF
C1043 gnd and2 0.08fF
C1044 comparator_0/fourinputOR_0/not_0/w_0_0# comparator_0/fourinputOR_0/not_0/in 0.06fF
C1045 vdd enableblock_0/enable1_0/AND_2/NAND_0/w_32_0# 0.05fF
C1046 comparator_0/AND_0/out comparator_0/XNOR_2/out 0.13fF
C1047 twotofourdecoder_0/AND_3/not_0/in OR_0/in1 0.02fF
C1048 gnd twotofourdecoder_0/AND_3/NAND_0/a_6_n14# 0.57fF
C1049 vdd twotofourdecoder_0/AND_2/not_0/w_0_0# 0.05fF
C1050 enableblock_2/enable1_1/AND_2/NAND_0/w_32_0# enableblock_2/enable1_1/AND_2/not_0/in 0.03fF
C1051 enableblock_1/enable1_1/AND_2/not_0/in comparator_0/A0 0.02fF
C1052 andblock_0/B3 enableblock_2/enable1_0/AND_1/not_0/in 0.02fF
C1053 vdd enableblock_0/enable1_1/AND_0/NAND_0/w_0_0# 0.05fF
C1054 addersubtractor_0/fulladder_2/AND_1/NAND_0/w_0_0# addersubtractor_0/fulladder_1/C 0.06fF
C1055 enableblock_2/enable1_1/AND_3/not_0/w_0_0# andblock_0/B0 0.03fF
C1056 vdd enableblock_1/enable1_0/AND_1/NAND_0/w_0_0# 0.05fF
C1057 gnd addersubtractor_0/XOR_1/NAND_0/a_6_n14# 0.57fF
C1058 vdd addersubtractor_0/fulladder_0/XOR_1/NAND_3/w_0_0# 0.05fF
C1059 gnd andblock_0/B0 0.28fF
C1060 vdd andblock_0/A3 0.26fF
C1061 addersubtractor_0/fulladder_0/XOR_0/NAND_3/w_0_0# vdd 0.05fF
C1062 addersubtractor_0/fulladder_0/XOR_1/in2 gnd 0.63fF
C1063 andblock_0/B0 andblock_0/AND_3/NAND_0/w_32_0# 0.06fF
C1064 andblock_0/B1 andblock_0/AND_2/NAND_0/w_32_0# 0.06fF
C1065 enableblock_0/enable1_1/AND_0/NAND_0/w_0_0# enableblock_0/enable1_1/AND_0/not_0/in 0.03fF
C1066 addersubtractor_0/fulladder_1/XOR_1/NAND_3/a_6_n14# gnd 0.57fF
C1067 enableblock_0/enable1_1/AND_2/not_0/w_0_0# enableblock_0/enable1_1/AND_2/not_0/in 0.06fF
C1068 enableblock_0/B_out3 addersubtractor_0/fulladder_2/XOR_0/NAND_1/w_0_0# 0.06fF
C1069 vdd addersubtractor_0/fulladder_1/XOR_1/NAND_3/w_32_0# 0.05fF
C1070 gnd XOR_0/NAND_3/in1 0.11fF
C1071 addersubtractor_0/fulladder_1/XOR_0/NAND_3/a_6_n14# gnd 0.57fF
C1072 vdd addersubtractor_0/fulladder_1/XOR_0/NAND_3/w_32_0# 0.05fF
C1073 vdd comparator_0/threeinputAND_0/not_0/w_0_0# 0.05fF
C1074 enableblock_0/A_out1 S0 0.06fF
C1075 vdd andblock_0/AND_3/not_0/in 0.29fF
C1076 gnd comparator_0/fourinputAND_1/fourinputNAND_0/a_6_n14# 0.47fF
C1077 addersubtractor_0/fulladder_0/AND_1/NAND_0/w_32_0# vdd 0.05fF
C1078 gnd enableblock_1/enable1_1/AND_1/not_0/in 0.04fF
C1079 addersubtractor_0/fulladder_2/XOR_1/NAND_3/w_32_0# addersubtractor_0/fulladder_2/XOR_1/NAND_3/in2 0.06fF
C1080 vdd OR_0/NOR_0/w_32_0# 0.03fF
C1081 A3 enableblock_2/enable1_0/AND_0/NAND_0/a_6_n14# 0.07fF
C1082 enableblock_0/enable1_0/AND_0/NAND_0/a_6_n14# enableblock_0/enable1_0/AND_0/not_0/in 0.12fF
C1083 B0 A2 0.19fF
C1084 gnd comparator_0/XNOR_0/XOR_0/NAND_2/in1 0.15fF
C1085 addersubtractor_0/fulladder_3/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_3/XOR_0/NAND_1/w_32_0# 0.06fF
C1086 vdd addersubtractor_0/fulladder_1/XOR_1/NAND_2/in1 0.25fF
C1087 comparator_0/fiveinputAND_0/fiveinputNAND_0/a_76_n14# comparator_0/XNOR_1/out 0.12fF
C1088 gnd comparator_0/fiveinputAND_0/not_0/in 0.01fF
C1089 addersubtractor_0/fulladder_2/XOR_1/NAND_0/a_6_n14# gnd 0.57fF
C1090 vdd comparator_0/fiveinputAND_0/fiveinputNAND_0/w_32_0# 0.05fF
C1091 gnd andblock_0/AND_1/NAND_0/a_6_n14# 0.57fF
C1092 adder2 addersubtractor_0/fulladder_2/XOR_1/NAND_3/a_6_n14# 0.12fF
C1093 addersubtractor_0/fulladder_2/XOR_0/NAND_3/w_32_0# addersubtractor_0/fulladder_2/XOR_0/NAND_3/in2 0.06fF
C1094 OR_0/out enableblock_0/enable1_1/AND_0/NAND_0/w_32_0# 0.06fF
C1095 vdd addersubtractor_0/fulladder_3/XOR_1/NAND_3/in2 0.25fF
C1096 comparator_0/A2 comparator_0/B2 2.42fF
C1097 comparator_0/fourinputAND_1/fourinputNAND_0/a_45_n14# comparator_0/XNOR_0/out 0.21fF
C1098 gnd enableblock_2/En 3.63fF
C1099 gnd addersubtractor_0/fulladder_3/XOR_1/NAND_2/in1 0.15fF
C1100 vdd addersubtractor_0/fulladder_3/XOR_0/NAND_3/in2 0.25fF
C1101 addersubtractor_0/fulladder_2/XOR_1/in2 addersubtractor_0/fulladder_2/XOR_0/NAND_3/a_6_n14# 0.12fF
C1102 comparator_0/threeinputAND_0/threeinputNAND_0/w_32_0# comparator_0/A2 0.06fF
C1103 enableblock_1/enable1_0/AND_1/NAND_0/w_0_0# enableblock_1/enable1_0/AND_1/not_0/in 0.03fF
C1104 vdd comparator_0/XNOR_1/XOR_0/NAND_3/in2 0.25fF
C1105 gnd comparator_0/fourinputAND_0/not_0/in 0.01fF
C1106 vdd comparator_0/not_2/out 0.07fF
C1107 vdd enableblock_0/enable1_1/AND_0/not_0/in 0.29fF
C1108 addersubtractor_0/fulladder_3/XOR_1/NAND_3/w_32_0# adder3 0.03fF
C1109 vdd addersubtractor_0/XOR_2/NAND_3/in2 0.25fF
C1110 twotofourdecoder_0/AND_3/NAND_0/a_6_n14# twotofourdecoder_0/AND_3/not_0/in 0.12fF
C1111 vdd addersubtractor_0/fulladder_2/XOR_1/NAND_0/w_0_0# 0.05fF
C1112 comparator_0/fourinputAND_0/fourinputNAND_0/w_100_0# comparator_0/XNOR_0/out 0.06fF
C1113 addersubtractor_0/fulladder_1/AND_0/not_0/w_0_0# addersubtractor_0/fulladder_1/AND_0/not_0/in 0.06fF
C1114 vdd comparator_0/XNOR_0/XOR_0/NAND_3/in2 0.25fF
C1115 addersubtractor_0/fulladder_3/XOR_0/NAND_3/w_32_0# addersubtractor_0/fulladder_3/XOR_1/in2 0.03fF
C1116 A1 B2 0.19fF
C1117 B0 A3 0.19fF
C1118 vdd andblock_0/B2 0.17fF
C1119 addersubtractor_0/XOR_0/NAND_0/w_0_0# enableblock_0/A_out2 0.06fF
C1120 gnd enableblock_0/enable1_0/AND_2/not_0/in 0.04fF
C1121 vdd XOR_0/in1 0.07fF
C1122 vdd XOR_0/NAND_1/w_0_0# 0.05fF
C1123 vdd comparator_0/XNOR_2/XOR_0/NAND_3/in2 0.25fF
C1124 AND_2/in2 AND_2/in1 0.06fF
C1125 enableblock_0/enable1_1/AND_1/NAND_0/w_32_0# enableblock_0/enable1_1/AND_1/not_0/in 0.03fF
C1126 addersubtractor_0/fulladder_0/C addersubtractor_0/fulladder_1/XOR_1/NAND_1/w_0_0# 0.06fF
C1127 gnd andblock_0/AND_1/not_0/in 0.04fF
C1128 comparator_0/XNOR_1/XOR_0/NAND_3/w_32_0# comparator_0/XNOR_1/not_0/in 0.03fF
C1129 comparator_0/fiveinputAND_0/not_0/in comparator_0/fiveinputAND_0/fiveinputNAND_0/w_100_0# 0.03fF
C1130 andblock_0/B3 andblock_0/A2 0.77fF
C1131 vdd comparator_0/XNOR_3/XOR_0/NAND_3/in2 0.25fF
C1132 vdd comparator_0/XNOR_0/XOR_0/NAND_1/w_32_0# 0.05fF
C1133 comparator_0/fourinputOR_0/in4 comparator_0/fiveinputAND_0/not_0/in 0.16fF
C1134 enableblock_2/enable1_0/AND_0/not_0/w_0_0# enableblock_2/enable1_0/AND_0/not_0/in 0.06fF
C1135 addersubtractor_0/XOR_2/NAND_1/w_0_0# enableblock_0/B_out2 0.06fF
C1136 enableblock_1/enable1_0/AND_0/NAND_0/w_32_0# enableblock_1/enable1_0/AND_0/not_0/in 0.03fF
C1137 addersubtractor_0/fulladder_0/AND_1/NAND_0/w_32_0# addersubtractor_0/fulladder_0/AND_1/not_0/in 0.03fF
C1138 vdd enableblock_0/enable1_1/AND_0/not_0/w_0_0# 0.05fF
C1139 vdd addersubtractor_0/XOR_3/NAND_1/w_0_0# 0.05fF
C1140 gnd comparator_0/XNOR_2/XOR_0/NAND_2/in1 0.15fF
C1141 enableblock_0/enable1_1/AND_1/not_0/w_0_0# enableblock_0/B_out2 0.03fF
C1142 vdd comparator_0/XNOR_2/XOR_0/NAND_1/w_32_0# 0.05fF
C1143 comparator_0/fourinputAND_1/fourinputNAND_0/w_32_0# comparator_0/XNOR_0/out 0.06fF
C1144 vdd enableblock_1/enable1_0/AND_1/not_0/in 0.29fF
C1145 S0 addersubtractor_0/XOR_3/NAND_0/w_32_0# 0.06fF
C1146 addersubtractor_0/fulladder_1/XOR_0/NAND_0/a_6_n14# gnd 0.57fF
C1147 addersubtractor_0/fulladder_0/AND_1/not_0/in vdd 0.29fF
C1148 vdd comparator_0/fourinputOR_0/fourinputNOR_0/a_45_6# 0.17fF
C1149 vdd addersubtractor_0/fulladder_1/AND_1/not_0/w_0_0# 0.05fF
C1150 gnd addersubtractor_0/fulladder_3/AND_0/NAND_0/a_6_n14# 0.57fF
C1151 vdd addersubtractor_0/fulladder_2/OR_0/in2 0.07fF
C1152 B2 S1 0.06fF
C1153 comparator_0/XNOR_0/XOR_0/NAND_3/w_32_0# comparator_0/XNOR_0/not_0/in 0.03fF
C1154 vdd comparator_0/XNOR_3/XOR_0/NAND_1/w_32_0# 0.05fF
C1155 addersubtractor_0/fulladder_2/XOR_1/NAND_1/w_0_0# addersubtractor_0/fulladder_2/XOR_1/NAND_3/in1 0.03fF
C1156 vdd comparator_0/XNOR_1/XOR_0/NAND_0/w_32_0# 0.05fF
C1157 vdd addersubtractor_0/fulladder_0/AND_0/not_0/in 0.03fF
C1158 AND_2/in2 comparator_0/A3 0.06fF
C1159 addersubtractor_0/fulladder_0/OR_0/NOR_0/w_0_0# vdd 0.05fF
C1160 gnd andblock_0/AND_2/NAND_0/a_6_n14# 0.57fF
C1161 vdd comparator_0/fourinputOR_0/not_0/in 0.10fF
C1162 vdd enableblock_2/enable1_1/AND_2/NAND_0/w_0_0# 0.05fF
C1163 enableblock_2/enable1_0/AND_3/not_0/w_0_0# enableblock_2/enable1_0/AND_3/not_0/in 0.06fF
C1164 addersubtractor_0/fulladder_2/AND_1/not_0/in gnd 0.04fF
C1165 enableblock_0/enable1_1/AND_0/not_0/w_0_0# enableblock_0/enable1_1/AND_0/not_0/in 0.06fF
C1166 addersubtractor_0/fulladder_2/XOR_0/NAND_1/w_0_0# addersubtractor_0/fulladder_2/XOR_0/NAND_3/in1 0.03fF
C1167 vdd comparator_0/fourinputAND_0/not_0/w_0_0# 0.05fF
C1168 vdd twotofourdecoder_0/AND_1/NAND_0/w_32_0# 0.05fF
C1169 B1 enableblock_2/En 0.13fF
C1170 A3 enableblock_0/enable1_1/AND_2/NAND_0/w_0_0# 0.06fF
C1171 vdd addersubtractor_0/fulladder_2/XOR_1/NAND_2/w_0_0# 0.05fF
C1172 comparator_0/XNOR_1/XOR_0/NAND_0/w_0_0# comparator_0/A2 0.06fF
C1173 XOR_0/NAND_1/w_0_0# XOR_0/in1 0.06fF
C1174 comparator_0/XNOR_2/XOR_0/NAND_3/w_32_0# comparator_0/XNOR_2/not_0/in 0.03fF
C1175 comparator_0/AND_0/not_0/w_0_0# comparator_0/AND_0/not_0/in 0.06fF
C1176 gnd enableblock_2/enable1_0/AND_0/NAND_0/a_6_n14# 0.57fF
C1177 OR_0/out A1 0.06fF
C1178 vdd enableblock_0/enable1_1/AND_3/not_0/w_0_0# 0.05fF
C1179 vdd enableblock_0/enable1_0/AND_0/NAND_0/w_0_0# 0.05fF
C1180 vdd addersubtractor_0/fulladder_2/XOR_0/NAND_2/w_0_0# 0.05fF
C1181 enableblock_2/En enableblock_2/enable1_1/AND_2/NAND_0/w_32_0# 0.06fF
C1182 vdd enableblock_0/B_out3 0.30fF
C1183 comparator_0/not_0/out comparator_0/B3 0.02fF
C1184 enableblock_0/enable1_1/AND_3/NAND_0/w_32_0# enableblock_0/enable1_1/AND_3/not_0/in 0.03fF
C1185 addersubtractor_0/XOR_2/NAND_1/a_6_n14# addersubtractor_0/XOR_2/NAND_3/in1 0.12fF
C1186 vdd addersubtractor_0/fulladder_3/XOR_0/NAND_2/in1 0.25fF
C1187 addersubtractor_0/fulladder_2/XOR_1/NAND_2/a_6_n14# addersubtractor_0/fulladder_2/XOR_1/NAND_3/in2 0.12fF
C1188 andblock_0/AND_2/not_0/in andblock_0/AND_2/NAND_0/w_32_0# 0.03fF
C1189 comparator_0/NOR_0/w_32_0# lesser 0.03fF
C1190 gnd addersubtractor_0/fulladder_3/XOR_1/NAND_2/a_6_n14# 0.59fF
C1191 vdd addersubtractor_0/fulladder_3/XOR_1/NAND_2/w_32_0# 0.05fF
C1192 comparator_0/not_3/out comparator_0/B0 0.02fF
C1193 enableblock_2/enable1_1/AND_1/NAND_0/a_6_n14# enableblock_2/enable1_1/AND_1/not_0/in 0.12fF
C1194 vdd addersubtractor_0/XOR_0/NAND_3/in1 0.25fF
C1195 gnd addersubtractor_0/fulladder_3/XOR_0/NAND_2/a_6_n14# 0.59fF
C1196 vdd addersubtractor_0/fulladder_2/OR_0/in1 0.12fF
C1197 comparator_0/XNOR_3/XOR_0/NAND_3/w_32_0# comparator_0/XNOR_3/not_0/in 0.03fF
C1198 vdd addersubtractor_0/fulladder_3/XOR_0/NAND_2/w_32_0# 0.05fF
C1199 addersubtractor_0/fulladder_2/XOR_0/NAND_2/a_6_n14# addersubtractor_0/fulladder_2/XOR_0/NAND_3/in2 0.12fF
C1200 vdd addersubtractor_0/fulladder_3/XOR_0/NAND_0/w_0_0# 0.05fF
C1201 addersubtractor_0/fulladder_2/AND_1/NAND_0/a_6_n14# addersubtractor_0/fulladder_2/AND_1/not_0/in 0.12fF
C1202 gnd comparator_0/XNOR_1/XOR_0/NAND_2/a_6_n14# 0.59fF
C1203 vdd comparator_0/XNOR_1/XOR_0/NAND_2/w_32_0# 0.05fF
C1204 gnd enableblock_2/enable1_0/AND_2/NAND_0/a_6_n14# 0.57fF
C1205 addersubtractor_0/fulladder_3/XOR_1/NAND_2/w_32_0# addersubtractor_0/fulladder_3/XOR_1/NAND_3/in2 0.03fF
C1206 addersubtractor_0/fulladder_3/OR_0/in2 addersubtractor_0/fulladder_3/OR_0/NOR_0/w_32_0# 0.06fF
C1207 vdd enableblock_2/enable1_0/AND_1/not_0/w_0_0# 0.05fF
C1208 enableblock_0/B_out3 enableblock_0/enable1_1/AND_0/not_0/in 0.02fF
C1209 gnd addersubtractor_0/XOR_2/NAND_2/a_6_n14# 0.59fF
C1210 vdd addersubtractor_0/XOR_2/NAND_2/w_32_0# 0.05fF
C1211 gnd comparator_0/XNOR_0/XOR_0/NAND_2/a_6_n14# 0.59fF
C1212 twotofourdecoder_0/AND_2/NAND_0/w_0_0# twotofourdecoder_0/AND_2/not_0/in 0.03fF
C1213 enableblock_0/A_out1 enableblock_0/enable1_0/AND_2/not_0/w_0_0# 0.03fF
C1214 addersubtractor_0/fulladder_1/AND_0/not_0/in addersubtractor_0/fulladder_1/AND_0/NAND_0/w_0_0# 0.03fF
C1215 vdd comparator_0/XNOR_0/XOR_0/NAND_2/w_32_0# 0.05fF
C1216 addersubtractor_0/XOR_2/out addersubtractor_0/XOR_2/NAND_3/w_32_0# 0.03fF
C1217 enableblock_1/enable1_1/AND_0/NAND_0/w_32_0# enableblock_1/enable1_1/AND_0/not_0/in 0.03fF
C1218 addersubtractor_0/fulladder_3/XOR_0/NAND_2/w_32_0# addersubtractor_0/fulladder_3/XOR_0/NAND_3/in2 0.03fF
C1219 enableblock_1/enable1_1/AND_3/not_0/w_0_0# enableblock_1/enable1_1/AND_3/not_0/in 0.06fF
C1220 gnd enableblock_1/enable1_1/AND_0/not_0/in 0.04fF
C1221 gnd twotofourdecoder_0/AND_0/not_0/in 0.04fF
C1222 addersubtractor_0/XOR_3/NAND_2/in1 addersubtractor_0/XOR_3/NAND_2/w_0_0# 0.06fF
C1223 gnd comparator_0/XNOR_2/XOR_0/NAND_2/a_6_n14# 0.59fF
C1224 gnd B0 0.76fF
C1225 vdd comparator_0/XNOR_2/XOR_0/NAND_2/w_32_0# 0.05fF
C1226 gnd AND_0/NAND_0/a_6_n14# 0.57fF
C1227 addersubtractor_0/fulladder_3/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_3/XOR_1/NAND_0/w_32_0# 0.03fF
C1228 vdd addersubtractor_0/XOR_1/NAND_3/w_0_0# 0.05fF
C1229 addersubtractor_0/XOR_0/out addersubtractor_0/fulladder_0/XOR_0/NAND_2/w_32_0# 0.06fF
C1230 comparator_0/XNOR_1/XOR_0/NAND_2/w_32_0# comparator_0/XNOR_1/XOR_0/NAND_3/in2 0.03fF
C1231 gnd comparator_0/XNOR_3/XOR_0/NAND_2/a_6_n14# 0.59fF
C1232 vdd comparator_0/XNOR_3/XOR_0/NAND_2/w_32_0# 0.05fF
C1233 gnd twotofourdecoder_0/AND_1/not_0/in 0.04fF
C1234 gnd enableblock_0/A_out0 0.82fF
C1235 addersubtractor_0/fulladder_1/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_1/XOR_0/NAND_0/a_6_n14# 0.12fF
C1236 addersubtractor_0/fulladder_1/AND_0/NAND_0/w_0_0# addersubtractor_0/XOR_1/out 0.06fF
C1237 S0 enableblock_0/A_out2 0.06fF
C1238 vdd comparator_0/AND_0/NAND_0/w_32_0# 0.05fF
C1239 addersubtractor_0/XOR_2/NAND_2/w_32_0# addersubtractor_0/XOR_2/NAND_3/in2 0.03fF
C1240 addersubtractor_0/fulladder_1/AND_0/NAND_0/w_32_0# enableblock_0/A_out1 0.06fF
C1241 enableblock_0/B_out3 enableblock_0/enable1_1/AND_0/not_0/w_0_0# 0.03fF
C1242 vdd addersubtractor_0/XOR_2/NAND_3/in1 0.29fF
C1243 AND_2/in2 comparator_0/AND_0/out 0.73fF
C1244 enableblock_2/enable1_0/AND_2/not_0/w_0_0# andblock_0/A2 0.03fF
C1245 addersubtractor_0/fulladder_1/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_1/XOR_1/NAND_3/w_0_0# 0.06fF
C1246 vdd enableblock_0/enable1_1/AND_1/NAND_0/w_32_0# 0.05fF
C1247 addersubtractor_0/fulladder_2/AND_0/not_0/in addersubtractor_0/fulladder_2/AND_0/NAND_0/w_32_0# 0.03fF
C1248 addersubtractor_0/fulladder_1/XOR_0/NAND_0/w_32_0# addersubtractor_0/XOR_1/out 0.06fF
C1249 addersubtractor_0/fulladder_0/OR_0/in2 addersubtractor_0/fulladder_0/OR_0/NOT_0/in 0.26fF
C1250 comparator_0/XNOR_0/XOR_0/NAND_2/w_32_0# comparator_0/XNOR_0/XOR_0/NAND_3/in2 0.03fF
C1251 enableblock_1/enable1_0/AND_2/not_0/w_0_0# comparator_0/A2 0.03fF
C1252 vdd AND_0/not_0/in 0.29fF
C1253 enableblock_2/enable1_1/AND_3/NAND_0/a_6_n14# enableblock_2/enable1_1/AND_3/not_0/in 0.12fF
C1254 comparator_0/XNOR_0/XOR_0/NAND_0/w_32_0# comparator_0/B3 0.06fF
C1255 addersubtractor_0/fulladder_1/XOR_0/NAND_3/in1 addersubtractor_0/fulladder_1/XOR_0/NAND_3/w_0_0# 0.06fF
C1256 addersubtractor_0/fulladder_1/AND_1/not_0/in addersubtractor_0/fulladder_1/OR_0/in1 0.02fF
C1257 addersubtractor_0/fulladder_3/AND_0/not_0/in addersubtractor_0/fulladder_3/OR_0/in2 0.02fF
C1258 A0 B2 0.19fF
C1259 vdd OR_0/in1 0.31fF
C1260 enableblock_0/enable1_0/AND_1/not_0/w_0_0# enableblock_0/enable1_0/AND_1/not_0/in 0.06fF
C1261 comparator_0/XNOR_2/XOR_0/NAND_2/w_32_0# comparator_0/XNOR_2/XOR_0/NAND_3/in2 0.03fF
C1262 vdd enableblock_2/enable1_1/AND_2/not_0/in 0.29fF
C1263 vdd addersubtractor_0/fulladder_1/OR_0/NOT_0/in 0.11fF
C1264 addersubtractor_0/fulladder_3/AND_1/NAND_0/w_0_0# addersubtractor_0/fulladder_3/AND_1/not_0/in 0.03fF
C1265 addersubtractor_0/fulladder_1/OR_0/NOR_0/w_0_0# addersubtractor_0/fulladder_1/OR_0/in1 0.06fF
C1266 addersubtractor_0/fulladder_1/C gnd 1.14fF
C1267 vdd enableblock_0/enable1_1/AND_2/NAND_0/w_32_0# 0.05fF
C1268 comparator_0/XNOR_2/XOR_0/NAND_0/w_32_0# comparator_0/B1 0.06fF
C1269 addersubtractor_0/XOR_0/NAND_2/in1 addersubtractor_0/XOR_0/NAND_0/a_6_n14# 0.12fF
C1270 vdd addersubtractor_0/fulladder_2/XOR_1/NAND_3/in1 0.25fF
C1271 vdd comparator_0/not_1/w_0_0# 0.05fF
C1272 vdd XOR_0/NAND_2/in1 0.25fF
C1273 gnd addersubtractor_0/fulladder_3/OR_0/NOT_0/in 0.60fF
C1274 vdd addersubtractor_0/fulladder_2/XOR_0/NAND_3/in1 0.25fF
C1275 addersubtractor_0/fulladder_0/C addersubtractor_0/fulladder_1/XOR_1/NAND_0/w_0_0# 0.06fF
C1276 comparator_0/XNOR_3/XOR_0/NAND_2/w_32_0# comparator_0/XNOR_3/XOR_0/NAND_3/in2 0.03fF
C1277 comparator_0/fourinputOR_0/fourinputNOR_0/a_13_6# comparator_0/fourinputOR_0/fourinputNOR_0/w_32_0# 0.03fF
C1278 addersubtractor_0/fulladder_2/OR_0/NOR_0/a_13_6# addersubtractor_0/fulladder_2/OR_0/NOR_0/w_0_0# 0.03fF
C1279 vdd enableblock_1/enable1_1/AND_1/NAND_0/w_0_0# 0.05fF
C1280 B0 B1 0.19fF
C1281 comparator_0/XNOR_3/XOR_0/NAND_0/w_32_0# comparator_0/B0 0.06fF
C1282 vdd comparator_0/not_0/w_0_0# 0.05fF
C1283 addersubtractor_0/fulladder_3/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_3/XOR_0/NAND_0/w_0_0# 0.03fF
C1284 AND_0/not_0/in XOR_0/in1 0.02fF
C1285 addersubtractor_0/XOR_1/NAND_0/w_32_0# S0 0.06fF
C1286 addersubtractor_0/fulladder_2/AND_1/NAND_0/a_6_n14# addersubtractor_0/fulladder_1/C 0.07fF
C1287 twotofourdecoder_0/not_0/out twotofourdecoder_0/AND_2/NAND_0/w_0_0# 0.06fF
C1288 enableblock_1/enable1_0/AND_2/NAND_0/w_0_0# A2 0.06fF
C1289 enableblock_0/B_out1 addersubtractor_0/XOR_3/out 0.11fF
C1290 vdd XOR_0/NAND_0/w_0_0# 0.05fF
C1291 addersubtractor_0/fulladder_3/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_3/XOR_1/NAND_1/w_32_0# 0.06fF
C1292 AND_0/in1 AND_0/NAND_0/w_0_0# 0.06fF
C1293 comparator_0/fourinputAND_1/fourinputNAND_0/w_63_0# comparator_0/XNOR_1/out 0.06fF
C1294 vdd enableblock_2/enable1_0/AND_3/NAND_0/w_32_0# 0.05fF
C1295 gnd enableblock_1/enable1_0/AND_1/NAND_0/a_6_n14# 0.57fF
C1296 vdd addersubtractor_0/XOR_2/NAND_2/in1 0.25fF
C1297 A2 B2 0.23fF
C1298 vdd enableblock_1/enable1_0/AND_0/not_0/w_0_0# 0.05fF
C1299 addersubtractor_0/fulladder_0/XOR_1/NAND_3/w_0_0# adder0 0.03fF
C1300 addersubtractor_0/fulladder_0/OR_0/NOT_0/in addersubtractor_0/fulladder_0/OR_0/NOT_0/w_0_0# 0.06fF
C1301 gnd OR_0/in2 0.34fF
C1302 vdd AND_2/NAND_0/w_0_0# 0.05fF
C1303 comparator_0/fourinputAND_1/not_0/in comparator_0/XNOR_1/out 0.03fF
C1304 S1 twotofourdecoder_0/not_1/out 0.16fF
C1305 vdd twotofourdecoder_0/AND_0/NAND_0/w_32_0# 0.05fF
C1306 addersubtractor_0/XOR_3/NAND_3/in1 addersubtractor_0/XOR_3/NAND_3/w_0_0# 0.06fF
C1307 vdd enableblock_0/enable1_0/AND_2/NAND_0/w_0_0# 0.05fF
C1308 addersubtractor_0/XOR_1/NAND_3/in1 addersubtractor_0/XOR_1/NAND_1/w_0_0# 0.03fF
C1309 vdd and2 0.18fF
C1310 addersubtractor_0/XOR_3/NAND_0/w_0_0# addersubtractor_0/XOR_3/NAND_2/in1 0.03fF
C1311 addersubtractor_0/fulladder_0/XOR_0/NAND_3/w_0_0# addersubtractor_0/fulladder_0/XOR_1/in2 0.03fF
C1312 enableblock_0/enable1_0/AND_0/NAND_0/w_32_0# enableblock_0/enable1_0/AND_0/not_0/in 0.03fF
C1313 enableblock_2/enable1_1/AND_2/NAND_0/w_0_0# enableblock_2/enable1_1/AND_2/not_0/in 0.03fF
C1314 XOR_0/NAND_3/w_32_0# Carry 0.03fF
C1315 S0 twotofourdecoder_0/not_0/out 0.02fF
C1316 andblock_0/AND_0/NAND_0/a_6_n14# andblock_0/AND_0/not_0/in 0.12fF
C1317 comparator_0/XNOR_2/not_0/w_0_0# comparator_0/XNOR_2/not_0/in 0.06fF
C1318 vdd comparator_0/not_3/w_0_0# 0.05fF
C1319 vdd enableblock_1/enable1_0/AND_3/not_0/w_0_0# 0.05fF
C1320 enableblock_1/enable1_0/AND_0/NAND_0/w_0_0# enableblock_1/enable1_0/AND_0/not_0/in 0.03fF
C1321 XOR_0/NAND_0/w_0_0# XOR_0/in1 0.06fF
C1322 addersubtractor_0/fulladder_0/AND_1/NAND_0/w_32_0# addersubtractor_0/fulladder_0/XOR_1/in2 0.06fF
C1323 vdd adder0 0.25fF
C1324 addersubtractor_0/fulladder_0/AND_0/not_0/w_0_0# addersubtractor_0/fulladder_0/AND_0/not_0/in 0.06fF
C1325 vdd andblock_0/B0 0.11fF
C1326 B2 A3 0.82fF
C1327 addersubtractor_0/fulladder_0/XOR_1/in2 vdd 0.47fF
C1328 addersubtractor_0/fulladder_3/AND_1/NAND_0/w_0_0# addersubtractor_0/fulladder_2/C 0.06fF
C1329 comparator_0/XNOR_3/not_0/w_0_0# comparator_0/XNOR_3/not_0/in 0.06fF
C1330 gnd comparator_0/fourinputOR_0/in2 0.16fF
C1331 gnd enableblock_0/enable1_1/AND_2/not_0/in 0.04fF
C1332 OR_0/out enableblock_0/enable1_0/AND_1/NAND_0/w_0_0# 0.06fF
C1333 enableblock_1/enable1_1/AND_3/not_0/in comparator_0/B0 0.02fF
C1334 vdd comparator_0/fourinputAND_1/fourinputNAND_0/w_100_0# 0.05fF
C1335 vdd addersubtractor_0/fulladder_2/XOR_1/NAND_3/w_0_0# 0.05fF
C1336 addersubtractor_0/fulladder_1/AND_1/NAND_0/a_6_n14# gnd 0.57fF
C1337 OR_0/out A2 0.07fF
C1338 enableblock_0/enable1_0/AND_2/NAND_0/w_32_0# enableblock_0/enable1_0/AND_2/not_0/in 0.03fF
C1339 gnd comparator_0/A2 1.18fF
C1340 vdd XOR_0/NAND_3/in1 0.25fF
C1341 vdd addersubtractor_0/fulladder_2/XOR_0/NAND_3/w_0_0# 0.05fF
C1342 addersubtractor_0/fulladder_2/XOR_1/in2 gnd 0.63fF
C1343 addersubtractor_0/fulladder_0/AND_1/NAND_0/w_0_0# vdd 0.05fF
C1344 comparator_0/NOR_0/a_13_6# lesser 0.04fF
C1345 enableblock_0/enable1_0/AND_3/not_0/w_0_0# enableblock_0/A_out0 0.03fF
C1346 vdd enableblock_1/enable1_1/AND_1/not_0/in 0.29fF
C1347 enableblock_0/enable1_0/AND_0/NAND_0/a_6_n14# A0 0.07fF
C1348 gnd addersubtractor_0/fulladder_3/XOR_1/NAND_3/a_6_n14# 0.57fF
C1349 comparator_0/threeinputAND_0/threeinputNAND_0/w_32_0# comparator_0/threeinputAND_0/not_0/in 0.03fF
C1350 vdd addersubtractor_0/fulladder_3/XOR_1/NAND_3/w_32_0# 0.05fF
C1351 enableblock_0/B_out1 addersubtractor_0/fulladder_3/XOR_0/NAND_1/w_0_0# 0.06fF
C1352 vdd comparator_0/XNOR_0/XOR_0/NAND_2/in1 0.25fF
C1353 vdd addersubtractor_0/fulladder_2/AND_1/NAND_0/w_32_0# 0.05fF
C1354 gnd addersubtractor_0/fulladder_3/XOR_0/NAND_3/a_6_n14# 0.57fF
C1355 vdd comparator_0/fiveinputAND_0/not_0/in 2.81fF
C1356 vdd addersubtractor_0/fulladder_3/XOR_0/NAND_3/w_32_0# 0.05fF
C1357 enableblock_0/B_out1 S0 0.06fF
C1358 comparator_0/XNOR_0/out comparator_0/B2 0.07fF
C1359 comparator_0/fiveinputAND_0/fiveinputNAND_0/w_32_0# comparator_0/fiveinputAND_0/not_0/in 0.03fF
C1360 gnd comparator_0/XNOR_1/XOR_0/NAND_3/a_6_n14# 0.57fF
C1361 addersubtractor_0/fulladder_3/XOR_1/NAND_3/w_32_0# addersubtractor_0/fulladder_3/XOR_1/NAND_3/in2 0.06fF
C1362 addersubtractor_0/fulladder_0/XOR_1/NAND_1/w_32_0# addersubtractor_0/fulladder_0/XOR_1/NAND_3/in1 0.03fF
C1363 OR_0/NOR_0/a_13_6# OR_0/NOT_0/in 0.04fF
C1364 vdd comparator_0/XNOR_1/XOR_0/NAND_3/w_32_0# 0.05fF
C1365 vdd comparator_0/fourinputAND_0/fourinputNAND_0/w_63_0# 0.05fF
C1366 gnd enableblock_2/enable1_1/AND_1/NAND_0/a_6_n14# 0.57fF
C1367 AND_0/in1 addersubtractor_0/fulladder_3/OR_0/NOT_0/in 0.02fF
C1368 addersubtractor_0/fulladder_1/AND_0/not_0/w_0_0# addersubtractor_0/fulladder_1/OR_0/in2 0.03fF
C1369 vdd enableblock_2/En 0.26fF
C1370 gnd addersubtractor_0/XOR_2/NAND_3/a_6_n14# 0.57fF
C1371 vdd addersubtractor_0/XOR_2/NAND_3/w_32_0# 0.05fF
C1372 addersubtractor_0/XOR_0/out addersubtractor_0/XOR_0/NAND_3/w_0_0# 0.03fF
C1373 comparator_0/fourinputOR_0/fourinputNOR_0/w_64_0# comparator_0/fourinputOR_0/fourinputNOR_0/a_77_6# 0.03fF
C1374 enableblock_1/enable1_0/AND_2/not_0/w_0_0# enableblock_1/enable1_0/AND_2/not_0/in 0.06fF
C1375 vdd addersubtractor_0/fulladder_3/XOR_1/NAND_2/in1 0.25fF
C1376 gnd comparator_0/XNOR_0/XOR_0/NAND_3/a_6_n14# 0.57fF
C1377 vdd comparator_0/XNOR_0/XOR_0/NAND_3/w_32_0# 0.05fF
C1378 B3 enableblock_2/En 0.13fF
C1379 addersubtractor_0/fulladder_3/XOR_0/NAND_3/w_32_0# addersubtractor_0/fulladder_3/XOR_0/NAND_3/in2 0.06fF
C1380 addersubtractor_0/fulladder_0/XOR_1/NAND_2/w_0_0# addersubtractor_0/fulladder_0/XOR_1/NAND_3/in2 0.03fF
C1381 addersubtractor_0/fulladder_0/XOR_0/NAND_1/w_32_0# addersubtractor_0/fulladder_0/XOR_0/NAND_3/in1 0.03fF
C1382 gnd enableblock_2/enable1_0/AND_3/not_0/in 0.04fF
C1383 OR_0/out A3 0.07fF
C1384 gnd comparator_0/B3 0.35fF
C1385 adder3 addersubtractor_0/fulladder_3/XOR_1/NAND_3/a_6_n14# 0.12fF
C1386 vdd comparator_0/fourinputAND_0/not_0/in 1.27fF
C1387 enableblock_1/enable1_1/AND_1/NAND_0/w_32_0# B1 0.06fF
C1388 addersubtractor_0/XOR_0/NAND_1/w_0_0# enableblock_0/A_out2 0.06fF
C1389 vdd AND_2/NAND_0/w_32_0# 0.05fF
C1390 vdd XOR_0/NAND_0/w_32_0# 0.05fF
C1391 gnd comparator_0/XNOR_2/XOR_0/NAND_3/a_6_n14# 0.57fF
C1392 vdd comparator_0/XNOR_2/XOR_0/NAND_3/w_32_0# 0.05fF
C1393 XOR_0/NAND_3/in1 XOR_0/NAND_1/w_0_0# 0.03fF
C1394 gnd comparator_0/B1 0.23fF
C1395 addersubtractor_0/fulladder_0/XOR_0/NAND_2/in1 gnd 0.15fF
C1396 addersubtractor_0/fulladder_0/XOR_0/NAND_2/w_0_0# addersubtractor_0/fulladder_0/XOR_0/NAND_3/in2 0.03fF
C1397 gnd andblock_0/AND_0/NAND_0/a_6_n14# 0.57fF
C1398 comparator_0/XNOR_1/XOR_0/NAND_3/w_32_0# comparator_0/XNOR_1/XOR_0/NAND_3/in2 0.06fF
C1399 addersubtractor_0/fulladder_3/XOR_1/in2 addersubtractor_0/fulladder_3/XOR_0/NAND_3/a_6_n14# 0.12fF
C1400 addersubtractor_0/fulladder_0/OR_0/NOT_0/in addersubtractor_0/fulladder_0/C 0.02fF
C1401 gnd comparator_0/XNOR_3/XOR_0/NAND_3/a_6_n14# 0.57fF
C1402 vdd comparator_0/fiveinputAND_0/fiveinputNAND_0/w_0_0# 0.05fF
C1403 comparator_0/fourinputAND_1/not_0/in comparator_0/XNOR_2/out 0.01fF
C1404 gnd addersubtractor_0/XOR_1/NAND_1/a_6_n14# 0.57fF
C1405 vdd comparator_0/XNOR_3/XOR_0/NAND_3/w_32_0# 0.05fF
C1406 XOR_0/NAND_2/w_32_0# XOR_0/NAND_3/in2 0.03fF
C1407 vdd twotofourdecoder_0/AND_1/NAND_0/w_0_0# 0.05fF
C1408 vdd enableblock_0/enable1_0/AND_2/not_0/in 0.29fF
C1409 gnd comparator_0/B0 0.22fF
C1410 addersubtractor_0/fulladder_1/AND_0/not_0/in gnd 0.04fF
C1411 addersubtractor_0/XOR_2/NAND_3/w_32_0# addersubtractor_0/XOR_2/NAND_3/in2 0.06fF
C1412 vdd enableblock_1/enable1_0/AND_2/NAND_0/w_32_0# 0.05fF
C1413 gnd enableblock_2/enable1_1/AND_2/NAND_0/a_6_n14# 0.57fF
C1414 addersubtractor_0/fulladder_2/AND_0/not_0/w_0_0# addersubtractor_0/fulladder_2/AND_0/not_0/in 0.06fF
C1415 addersubtractor_0/fulladder_0/XOR_0/NAND_0/w_32_0# vdd 0.05fF
C1416 comparator_0/XNOR_1/not_0/in comparator_0/XNOR_1/XOR_0/NAND_3/a_6_n14# 0.12fF
C1417 vdd twotofourdecoder_0/not_1/w_0_0# 0.05fF
C1418 vdd enableblock_2/enable1_1/AND_1/not_0/w_0_0# 0.05fF
C1419 vdd andblock_0/AND_1/not_0/in 0.29fF
C1420 comparator_0/XNOR_0/XOR_0/NAND_2/in1 comparator_0/XNOR_0/XOR_0/NAND_1/w_32_0# 0.06fF
C1421 vdd comparator_0/fourinputAND_1/fourinputNAND_0/w_0_0# 0.05fF
C1422 enableblock_2/enable1_0/AND_2/NAND_0/a_6_n14# enableblock_2/enable1_0/AND_2/not_0/in 0.12fF
C1423 addersubtractor_0/fulladder_0/AND_1/NAND_0/w_0_0# addersubtractor_0/fulladder_0/AND_1/not_0/in 0.03fF
C1424 comparator_0/XNOR_0/XOR_0/NAND_3/w_32_0# comparator_0/XNOR_0/XOR_0/NAND_3/in2 0.06fF
C1425 S0 twotofourdecoder_0/AND_0/NAND_0/w_0_0# 0.06fF
C1426 vdd addersubtractor_0/fulladder_0/XOR_1/NAND_0/w_32_0# 0.05fF
C1427 vdd XOR_0/NAND_2/w_0_0# 0.05fF
C1428 vdd comparator_0/XNOR_2/XOR_0/NAND_2/in1 0.25fF
C1429 vdd enableblock_1/enable1_1/AND_0/NAND_0/w_0_0# 0.05fF
C1430 enableblock_1/enable1_0/AND_0/not_0/in comparator_0/A3 0.02fF
C1431 gnd greater 0.08fF
C1432 addersubtractor_0/fulladder_1/C addersubtractor_0/fulladder_2/XOR_1/NAND_1/w_0_0# 0.06fF
C1433 addersubtractor_0/XOR_1/out gnd 0.56fF
C1434 vdd twotofourdecoder_0/not_0/w_0_0# 0.05fF
C1435 addersubtractor_0/fulladder_1/AND_1/NAND_0/w_32_0# addersubtractor_0/fulladder_1/AND_1/not_0/in 0.03fF
C1436 gnd B2 0.83fF
C1437 addersubtractor_0/fulladder_0/AND_1/not_0/w_0_0# addersubtractor_0/fulladder_0/OR_0/in1 0.03fF
C1438 vdd vdd 0.05fF
C1439 comparator_0/XNOR_0/not_0/in comparator_0/XNOR_0/XOR_0/NAND_3/a_6_n14# 0.12fF
C1440 gnd comparator_0/fourinputOR_0/in3 0.79fF
C1441 vdd addersubtractor_0/fulladder_2/AND_0/NAND_0/w_32_0# 0.05fF
C1442 comparator_0/XNOR_2/XOR_0/NAND_3/w_32_0# comparator_0/XNOR_2/XOR_0/NAND_3/in2 0.06fF
C1443 gnd enableblock_0/B_out0 0.82fF
C1444 addersubtractor_0/XOR_0/NAND_2/in1 gnd 0.15fF
C1445 vdd addersubtractor_0/fulladder_1/OR_0/NOT_0/w_0_0# 0.05fF
C1446 AND_2/in1 comparator_0/fourinputAND_1/not_0/in 0.02fF
C1447 vdd addersubtractor_0/fulladder_2/AND_1/not_0/in 0.29fF
C1448 S0 enableblock_0/B_out2 0.06fF
C1449 gnd addersubtractor_0/fulladder_3/XOR_0/NAND_0/a_6_n14# 0.57fF
C1450 vdd addersubtractor_0/fulladder_3/AND_1/not_0/w_0_0# 0.05fF
C1451 enableblock_1/enable1_1/AND_2/NAND_0/w_0_0# A0 0.06fF
C1452 addersubtractor_0/fulladder_3/XOR_1/NAND_1/w_0_0# addersubtractor_0/fulladder_3/XOR_1/NAND_3/in1 0.03fF
C1453 comparator_0/XNOR_2/not_0/in comparator_0/XNOR_2/XOR_0/NAND_3/a_6_n14# 0.12fF
C1454 AND_2/in2 twotofourdecoder_0/AND_1/not_0/w_0_0# 0.03fF
C1455 vdd addersubtractor_0/fulladder_2/OR_0/NOR_0/w_0_0# 0.05fF
C1456 andblock_0/AND_0/NAND_0/w_32_0# andblock_0/AND_0/not_0/in 0.03fF
C1457 comparator_0/XNOR_3/XOR_0/NAND_3/w_32_0# comparator_0/XNOR_3/XOR_0/NAND_3/in2 0.06fF
C1458 enableblock_0/enable1_1/AND_3/NAND_0/w_0_0# enableblock_0/enable1_1/AND_3/not_0/in 0.03fF
C1459 enableblock_0/enable1_0/AND_3/NAND_0/w_32_0# B1 0.06fF
C1460 vdd AND_0/NAND_0/w_0_0# 0.05fF
C1461 addersubtractor_0/fulladder_3/XOR_0/NAND_1/w_0_0# addersubtractor_0/fulladder_3/XOR_0/NAND_3/in1 0.03fF
C1462 gnd andblock_0/B3 0.44fF
C1463 addersubtractor_0/XOR_0/NAND_2/in1 addersubtractor_0/XOR_0/NAND_1/w_32_0# 0.06fF
C1464 equal AND_2/not_0/in 0.02fF
C1465 enableblock_1/enable1_1/AND_2/NAND_0/a_6_n14# enableblock_1/enable1_1/AND_2/not_0/in 0.12fF
C1466 comparator_0/XNOR_0/not_0/w_0_0# comparator_0/XNOR_0/not_0/in 0.06fF
C1467 addersubtractor_0/XOR_1/NAND_0/w_32_0# addersubtractor_0/XOR_1/NAND_2/in1 0.03fF
C1468 comparator_0/XNOR_3/not_0/in comparator_0/XNOR_3/XOR_0/NAND_3/a_6_n14# 0.12fF
C1469 XOR_0/NAND_2/in1 XOR_0/NAND_0/w_0_0# 0.03fF
C1470 comparator_0/fourinputAND_0/not_0/w_0_0# comparator_0/fourinputAND_0/not_0/in 0.06fF
C1471 addersubtractor_0/fulladder_0/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_0/XOR_0/NAND_2/w_0_0# 0.06fF
C1472 comparator_0/XNOR_1/XOR_0/NAND_2/in1 comparator_0/XNOR_1/XOR_0/NAND_2/w_0_0# 0.06fF
C1473 comparator_0/XNOR_1/XOR_0/NAND_1/w_0_0# comparator_0/XNOR_1/XOR_0/NAND_3/in1 0.03fF
C1474 enableblock_1/enable1_1/AND_0/NAND_0/a_6_n14# enableblock_1/enable1_1/AND_0/not_0/in 0.12fF
C1475 addersubtractor_0/fulladder_3/XOR_1/NAND_2/a_6_n14# addersubtractor_0/fulladder_3/XOR_1/NAND_3/in2 0.12fF
C1476 twotofourdecoder_0/AND_3/not_0/w_0_0# twotofourdecoder_0/AND_3/not_0/in 0.06fF
C1477 twotofourdecoder_0/AND_0/NAND_0/a_6_n14# twotofourdecoder_0/AND_0/not_0/in 0.12fF
C1478 gnd OR_0/out 3.60fF
C1479 comparator_0/XNOR_2/XOR_0/NAND_2/in1 comparator_0/XNOR_2/XOR_0/NAND_1/w_32_0# 0.06fF
C1480 AND_2/in2 enableblock_1/enable1_0/AND_3/NAND_0/w_0_0# 0.06fF
C1481 comparator_0/B2 comparator_0/A1 0.76fF
C1482 addersubtractor_0/XOR_2/out addersubtractor_0/XOR_2/NAND_3/a_6_n14# 0.12fF
C1483 AND_2/in1 comparator_0/fourinputAND_1/not_0/w_0_0# 0.03fF
C1484 addersubtractor_0/fulladder_3/XOR_0/NAND_2/a_6_n14# addersubtractor_0/fulladder_3/XOR_0/NAND_3/in2 0.12fF
C1485 addersubtractor_0/fulladder_3/AND_1/NAND_0/a_6_n14# addersubtractor_0/fulladder_3/AND_1/not_0/in 0.12fF
C1486 andblock_0/B1 enableblock_2/enable1_1/AND_1/not_0/in 0.02fF
C1487 enableblock_0/A_out3 addersubtractor_0/fulladder_0/XOR_0/NAND_0/w_0_0# 0.06fF
C1488 vdd enableblock_1/enable1_1/AND_0/not_0/in 0.29fF
C1489 vdd twotofourdecoder_0/AND_0/not_0/in 0.29fF
C1490 enableblock_1/enable1_0/AND_3/NAND_0/w_32_0# enableblock_1/enable1_0/AND_3/not_0/in 0.03fF
C1491 comparator_0/fourinputAND_0/fourinputNAND_0/w_32_0# comparator_0/A1 0.06fF
C1492 B0 B3 0.19fF
C1493 B1 B2 0.19fF
C1494 comparator_0/XNOR_1/XOR_0/NAND_2/a_6_n14# comparator_0/XNOR_1/XOR_0/NAND_3/in2 0.12fF
C1495 comparator_0/fourinputOR_0/fourinputNOR_0/w_64_0# comparator_0/fourinputOR_0/in3 0.06fF
C1496 addersubtractor_0/fulladder_2/AND_0/not_0/in addersubtractor_0/fulladder_2/AND_0/NAND_0/w_0_0# 0.03fF
C1497 vdd twotofourdecoder_0/AND_1/not_0/in 0.29fF
C1498 enableblock_2/enable1_0/AND_1/NAND_0/w_0_0# enableblock_2/enable1_0/AND_1/not_0/in 0.03fF
C1499 vdd enableblock_0/A_out0 0.17fF
C1500 addersubtractor_0/fulladder_0/XOR_1/NAND_1/a_6_n14# gnd 0.57fF
C1501 vdd addersubtractor_0/fulladder_0/XOR_1/NAND_1/w_32_0# 0.05fF
C1502 S0 A1 0.16fF
C1503 gnd enableblock_1/enable1_0/AND_2/not_0/in 0.04fF
C1504 addersubtractor_0/XOR_3/NAND_1/w_32_0# addersubtractor_0/XOR_3/NAND_3/in1 0.03fF
C1505 addersubtractor_0/XOR_2/NAND_2/a_6_n14# addersubtractor_0/XOR_2/NAND_3/in2 0.12fF
C1506 addersubtractor_0/fulladder_0/OR_0/NOT_0/in addersubtractor_0/fulladder_0/OR_0/NOR_0/w_32_0# 0.03fF
C1507 addersubtractor_0/fulladder_0/XOR_0/NAND_1/a_6_n14# gnd 0.57fF
C1508 addersubtractor_0/fulladder_0/XOR_0/NAND_1/w_32_0# vdd 0.05fF
C1509 S0 twotofourdecoder_0/AND_3/NAND_0/w_32_0# 0.06fF
C1510 addersubtractor_0/XOR_1/out addersubtractor_0/fulladder_1/XOR_0/NAND_2/w_32_0# 0.06fF
C1511 comparator_0/XNOR_0/XOR_0/NAND_2/a_6_n14# comparator_0/XNOR_0/XOR_0/NAND_3/in2 0.12fF
C1512 addersubtractor_0/XOR_3/NAND_2/in1 addersubtractor_0/XOR_3/NAND_0/a_6_n14# 0.12fF
C1513 addersubtractor_0/fulladder_2/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_2/XOR_0/NAND_0/a_6_n14# 0.12fF
C1514 addersubtractor_0/fulladder_2/AND_0/NAND_0/w_0_0# addersubtractor_0/XOR_2/out 0.06fF
C1515 vdd enableblock_1/enable1_1/AND_0/not_0/w_0_0# 0.05fF
C1516 vdd enableblock_2/enable1_1/AND_3/NAND_0/w_32_0# 0.05fF
C1517 addersubtractor_0/fulladder_2/AND_0/NAND_0/w_32_0# enableblock_0/B_out3 0.06fF
C1518 addersubtractor_0/fulladder_2/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_2/XOR_1/NAND_3/w_0_0# 0.06fF
C1519 addersubtractor_0/fulladder_3/AND_0/not_0/in addersubtractor_0/fulladder_3/AND_0/NAND_0/w_32_0# 0.03fF
C1520 addersubtractor_0/fulladder_2/XOR_0/NAND_0/w_32_0# addersubtractor_0/XOR_2/out 0.06fF
C1521 vdd comparator_0/AND_0/not_0/w_0_0# 0.05fF
C1522 comparator_0/XNOR_2/XOR_0/NAND_2/a_6_n14# comparator_0/XNOR_2/XOR_0/NAND_3/in2 0.12fF
C1523 comparator_0/XNOR_3/XOR_0/NAND_2/in1 comparator_0/XNOR_3/XOR_0/NAND_0/w_0_0# 0.03fF
C1524 comparator_0/fiveinputAND_0/fiveinputNAND_0/a_6_n14# comparator_0/A0 0.04fF
C1525 vdd addersubtractor_0/fulladder_1/C 0.18fF
C1526 vdd enableblock_0/enable1_1/AND_2/NAND_0/w_0_0# 0.05fF
C1527 addersubtractor_0/fulladder_2/XOR_0/NAND_3/in1 addersubtractor_0/fulladder_2/XOR_0/NAND_3/w_0_0# 0.06fF
C1528 addersubtractor_0/fulladder_2/AND_1/not_0/in addersubtractor_0/fulladder_2/OR_0/in1 0.02fF
C1529 comparator_0/not_0/out comparator_0/AND_0/NAND_0/w_0_0# 0.06fF
C1530 vdd enableblock_2/enable1_0/AND_1/NAND_0/w_32_0# 0.05fF
C1531 OR_0/out B1 0.07fF
C1532 vdd addersubtractor_0/XOR_0/NAND_2/w_0_0# 0.05fF
C1533 twotofourdecoder_0/AND_2/not_0/w_0_0# OR_0/in2 0.03fF
C1534 gnd enableblock_0/enable1_0/AND_0/NAND_0/a_6_n14# 0.57fF
C1535 AND_2/in2 A1 0.06fF
C1536 enableblock_1/enable1_0/AND_0/NAND_0/w_0_0# A3 0.06fF
C1537 comparator_0/XNOR_3/XOR_0/NAND_2/a_6_n14# comparator_0/XNOR_3/XOR_0/NAND_3/in2 0.12fF
C1538 B3 enableblock_2/enable1_0/AND_1/NAND_0/w_32_0# 0.06fF
C1539 vdd enableblock_1/enable1_1/AND_3/not_0/w_0_0# 0.05fF
C1540 enableblock_1/enable1_1/AND_1/NAND_0/w_0_0# enableblock_1/enable1_1/AND_1/not_0/in 0.03fF
C1541 vdd addersubtractor_0/fulladder_3/OR_0/NOT_0/in 0.11fF
C1542 addersubtractor_0/fulladder_2/OR_0/NOR_0/w_0_0# addersubtractor_0/fulladder_2/OR_0/in1 0.06fF
C1543 enableblock_0/enable1_0/AND_3/NAND_0/a_6_n14# enableblock_0/enable1_0/AND_3/not_0/in 0.12fF
C1544 S0 addersubtractor_0/XOR_3/NAND_2/w_32_0# 0.06fF
C1545 vdd comparator_0/XNOR_2/not_0/w_0_0# 0.05fF
C1546 XOR_0/NAND_0/w_32_0# OR_0/in1 0.06fF
C1547 OR_0/out OR_0/NOT_0/w_0_0# 0.03fF
C1548 addersubtractor_0/fulladder_1/C addersubtractor_0/fulladder_2/XOR_1/NAND_0/w_0_0# 0.06fF
C1549 vdd comparator_0/XNOR_3/not_0/w_0_0# 0.05fF
C1550 addersubtractor_0/XOR_0/NAND_2/w_32_0# S0 0.06fF
C1551 addersubtractor_0/fulladder_3/OR_0/NOR_0/a_13_6# addersubtractor_0/fulladder_3/OR_0/NOR_0/w_0_0# 0.03fF
C1552 and1 andblock_0/AND_2/not_0/in 0.02fF
C1553 OR_0/out enableblock_0/enable1_1/AND_1/NAND_0/w_0_0# 0.06fF
C1554 AND_0/in1 addersubtractor_0/fulladder_3/OR_0/NOT_0/w_0_0# 0.03fF
C1555 gnd enableblock_0/enable1_0/AND_2/NAND_0/a_6_n14# 0.57fF
C1556 andblock_0/AND_0/not_0/w_0_0# andblock_0/AND_0/not_0/in 0.06fF
C1557 gnd comparator_0/XNOR_1/out 0.69fF
C1558 twotofourdecoder_0/not_1/out twotofourdecoder_0/AND_3/NAND_0/w_0_0# 0.06fF
C1559 vdd enableblock_0/enable1_0/AND_1/not_0/w_0_0# 0.05fF
C1560 vdd comparator_0/NOR_0/w_0_0# 0.05fF
C1561 enableblock_2/enable1_0/AND_0/not_0/in enableblock_2/enable1_0/AND_0/NAND_0/w_0_0# 0.03fF
C1562 XOR_0/NAND_2/in1 XOR_0/NAND_0/w_32_0# 0.03fF
C1563 addersubtractor_0/fulladder_0/OR_0/NOT_0/in addersubtractor_0/fulladder_0/OR_0/NOR_0/a_13_6# 0.04fF
C1564 addersubtractor_0/fulladder_3/AND_1/NAND_0/a_6_n14# addersubtractor_0/fulladder_2/C 0.07fF
C1565 AND_2/in1 lesser 0.13fF
C1566 twotofourdecoder_0/AND_1/NAND_0/w_32_0# twotofourdecoder_0/AND_1/not_0/in 0.03fF
C1567 vdd enableblock_2/enable1_0/AND_3/NAND_0/w_0_0# 0.05fF
C1568 vdd comparator_0/NOR_0/w_32_0# 0.03fF
C1569 comparator_0/fourinputOR_0/not_0/w_0_0# greater 0.03fF
C1570 gnd enableblock_2/enable1_0/AND_0/not_0/in 0.04fF
C1571 andblock_0/A1 enableblock_2/enable1_1/AND_0/not_0/in 0.02fF
C1572 addersubtractor_0/XOR_3/NAND_1/w_32_0# addersubtractor_0/XOR_3/NAND_2/in1 0.06fF
C1573 OR_0/in2 OR_0/NOR_0/w_32_0# 0.06fF
C1574 gnd twotofourdecoder_0/not_1/out 3.35fF
C1575 gnd addersubtractor_0/XOR_1/NAND_3/in1 0.11fF
C1576 addersubtractor_0/fulladder_0/OR_0/NOT_0/w_0_0# addersubtractor_0/fulladder_0/C 0.03fF
C1577 vdd OR_0/in2 0.33fF
C1578 XOR_0/NAND_3/w_32_0# XOR_0/NAND_3/in2 0.06fF
C1579 enableblock_2/enable1_1/AND_0/NAND_0/w_32_0# enableblock_2/enable1_1/AND_0/not_0/in 0.03fF
C1580 enableblock_2/enable1_1/AND_3/not_0/w_0_0# enableblock_2/enable1_1/AND_3/not_0/in 0.06fF
C1581 enableblock_0/enable1_0/AND_1/NAND_0/w_32_0# enableblock_0/enable1_0/AND_1/not_0/in 0.03fF
C1582 XOR_0/NAND_2/in1 XOR_0/NAND_2/w_0_0# 0.06fF
C1583 addersubtractor_0/fulladder_1/XOR_1/NAND_3/w_0_0# adder1 0.03fF
C1584 addersubtractor_0/fulladder_1/OR_0/NOT_0/in addersubtractor_0/fulladder_1/OR_0/NOT_0/w_0_0# 0.06fF
C1585 vdd comparator_0/fourinputOR_0/fourinputNOR_0/a_77_6# 0.18fF
C1586 Carry XOR_0/NAND_3/a_6_n14# 0.12fF
C1587 vdd addersubtractor_0/fulladder_0/XOR_1/NAND_3/in2 0.25fF
C1588 vdd XOR_0/NAND_3/w_0_0# 0.05fF
C1589 comparator_0/XNOR_1/not_0/in comparator_0/XNOR_1/out 0.02fF
C1590 vdd enableblock_1/enable1_1/AND_1/NAND_0/w_32_0# 0.05fF
C1591 gnd enableblock_2/enable1_1/AND_3/not_0/in 0.04fF
C1592 AND_0/not_0/in AND_0/NAND_0/w_0_0# 0.03fF
C1593 addersubtractor_0/fulladder_0/XOR_1/NAND_2/in1 gnd 0.15fF
C1594 addersubtractor_0/fulladder_0/XOR_0/NAND_3/in2 vdd 0.25fF
C1595 gnd comparator_0/threeinputAND_0/not_0/in 0.75fF
C1596 addersubtractor_0/XOR_3/NAND_0/w_32_0# addersubtractor_0/XOR_3/NAND_2/in1 0.03fF
C1597 vdd addersubtractor_0/fulladder_2/AND_0/not_0/w_0_0# 0.05fF
C1598 addersubtractor_0/fulladder_1/XOR_0/NAND_3/w_0_0# addersubtractor_0/fulladder_1/XOR_1/in2 0.03fF
C1599 enableblock_2/enable1_1/AND_0/not_0/w_0_0# andblock_0/A1 0.03fF
C1600 addersubtractor_0/fulladder_0/AND_1/NAND_0/a_6_n14# gnd 0.57fF
C1601 addersubtractor_0/fulladder_0/OR_0/in2 addersubtractor_0/fulladder_0/OR_0/NOR_0/w_32_0# 0.06fF
C1602 addersubtractor_0/fulladder_0/AND_0/not_0/w_0_0# vdd 0.05fF
C1603 comparator_0/threeinputAND_0/not_0/w_0_0# comparator_0/fourinputOR_0/in2 0.03fF
C1604 andblock_0/A2 andblock_0/AND_1/NAND_0/w_0_0# 0.06fF
C1605 addersubtractor_0/fulladder_0/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_0/XOR_1/NAND_0/w_0_0# 0.03fF
C1606 addersubtractor_0/fulladder_1/AND_1/NAND_0/w_32_0# addersubtractor_0/fulladder_1/XOR_1/in2 0.06fF
C1607 S0 A0 0.13fF
C1608 vdd comparator_0/fourinputOR_0/in2 0.95fF
C1609 gnd comparator_0/XNOR_0/out 0.98fF
C1610 vdd enableblock_0/enable1_1/AND_2/not_0/in 0.29fF
C1611 addersubtractor_0/fulladder_0/AND_1/not_0/w_0_0# vdd 0.05fF
C1612 A1 enableblock_2/enable1_1/AND_0/NAND_0/a_6_n14# 0.07fF
C1613 vdd enableblock_1/enable1_1/AND_2/NAND_0/w_32_0# 0.05fF
C1614 vdd addersubtractor_0/XOR_3/NAND_2/w_0_0# 0.05fF
C1615 vdd adder2 0.25fF
C1616 enableblock_0/enable1_0/AND_2/NAND_0/w_0_0# enableblock_0/enable1_0/AND_2/not_0/in 0.03fF
C1617 vdd comparator_0/A2 0.20fF
C1618 vdd addersubtractor_0/fulladder_1/OR_0/NOR_0/w_32_0# 0.03fF
C1619 vdd addersubtractor_0/fulladder_2/XOR_1/in2 0.47fF
C1620 vdd comparator_0/threeinputAND_0/threeinputNAND_0/w_0_0# 0.05fF
C1621 enableblock_1/enable1_0/AND_1/NAND_0/a_6_n14# enableblock_1/enable1_0/AND_1/not_0/in 0.12fF
C1622 AND_0/NAND_0/a_6_n14# AND_0/not_0/in 0.12fF
C1623 andblock_0/AND_1/not_0/in and2 0.02fF
C1624 vdd comparator_0/fourinputAND_0/fourinputNAND_0/w_0_0# 0.05fF
C1625 gnd addersubtractor_0/XOR_0/NAND_1/a_6_n14# 0.57fF
C1626 addersubtractor_0/fulladder_3/AND_1/NAND_0/a_6_n14# gnd 0.57fF
C1627 comparator_0/XNOR_1/not_0/w_0_0# comparator_0/XNOR_1/out 0.03fF
C1628 addersubtractor_0/XOR_3/out addersubtractor_0/XOR_3/NAND_3/w_32_0# 0.03fF
C1629 vdd comparator_0/threeinputAND_0/threeinputNAND_0/w_63_0# 0.05fF
C1630 comparator_0/not_1/out comparator_0/B2 0.02fF
C1631 andblock_0/A3 andblock_0/AND_0/NAND_0/a_6_n14# 0.07fF
C1632 gnd comparator_0/fourinputAND_0/fourinputNAND_0/a_76_n14# 0.04fF
C1633 gnd andblock_0/A1 0.22fF
C1634 addersubtractor_0/fulladder_0/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_0/XOR_1/NAND_1/a_6_n14# 0.12fF
C1635 vdd addersubtractor_0/XOR_1/NAND_0/w_0_0# 0.05fF
C1636 S1 twotofourdecoder_0/not_0/out 0.14fF
C1637 gnd addersubtractor_0/XOR_3/NAND_0/a_6_n14# 0.57fF
C1638 andblock_0/AND_0/not_0/w_0_0# and3 0.03fF
C1639 comparator_0/fourinputOR_0/fourinputNOR_0/a_77_6# comparator_0/fourinputOR_0/fourinputNOR_0/a_45_6# 0.04fF
C1640 vdd comparator_0/fiveinputAND_0/fiveinputNAND_0/w_133_0# 0.05fF
C1641 gnd comparator_0/XNOR_2/out 0.31fF
C1642 enableblock_2/enable1_1/AND_2/not_0/w_0_0# andblock_0/A0 0.03fF
C1643 addersubtractor_0/fulladder_1/OR_0/in2 gnd 0.36fF
C1644 addersubtractor_0/fulladder_0/XOR_0/NAND_3/in1 addersubtractor_0/fulladder_0/XOR_0/NAND_1/a_6_n14# 0.12fF
C1645 comparator_0/fourinputAND_0/fourinputNAND_0/w_0_0# comparator_0/not_2/out 0.06fF
C1646 vdd enableblock_2/enable1_0/AND_3/not_0/in 0.29fF
C1647 AND_2/in2 A0 0.06fF
C1648 vdd comparator_0/B3 0.26fF
C1649 comparator_0/XNOR_0/out comparator_0/fiveinputAND_0/fiveinputNAND_0/w_100_0# 0.06fF
C1650 addersubtractor_0/fulladder_1/XOR_1/NAND_1/w_32_0# addersubtractor_0/fulladder_1/XOR_1/NAND_3/in1 0.03fF
C1651 comparator_0/XNOR_0/out comparator_0/XNOR_0/not_0/in 0.02fF
C1652 comparator_0/fourinputOR_0/fourinputNOR_0/a_77_6# comparator_0/fourinputOR_0/not_0/in 0.04fF
C1653 vdd enableblock_0/enable1_0/AND_3/NAND_0/w_32_0# 0.05fF
C1654 addersubtractor_0/fulladder_2/AND_0/not_0/w_0_0# addersubtractor_0/fulladder_2/OR_0/in2 0.03fF
C1655 addersubtractor_0/fulladder_0/XOR_1/NAND_2/in1 addersubtractor_0/fulladder_0/XOR_1/NAND_2/w_0_0# 0.06fF
C1656 comparator_0/AND_0/NAND_0/a_6_n14# comparator_0/AND_0/not_0/in 0.12fF
C1657 addersubtractor_0/fulladder_0/XOR_1/in2 addersubtractor_0/fulladder_0/XOR_1/NAND_0/w_32_0# 0.06fF
C1658 andblock_0/AND_0/NAND_0/w_0_0# andblock_0/AND_0/not_0/in 0.03fF
C1659 comparator_0/fourinputAND_1/fourinputNAND_0/w_32_0# comparator_0/fourinputAND_1/not_0/in 0.03fF
C1660 comparator_0/AND_0/NAND_0/w_0_0# comparator_0/AND_0/not_0/in 0.03fF
C1661 gnd andblock_0/B1 0.38fF
C1662 vdd comparator_0/B1 0.35fF
C1663 addersubtractor_0/XOR_1/NAND_1/w_32_0# addersubtractor_0/XOR_1/NAND_3/in1 0.03fF
C1664 addersubtractor_0/fulladder_0/XOR_0/NAND_2/in1 vdd 0.25fF
C1665 comparator_0/fourinputAND_0/fourinputNAND_0/w_63_0# comparator_0/fourinputAND_0/not_0/in 0.03fF
C1666 vdd twotofourdecoder_0/AND_3/not_0/w_0_0# 0.05fF
C1667 addersubtractor_0/fulladder_1/XOR_1/NAND_2/w_0_0# addersubtractor_0/fulladder_1/XOR_1/NAND_3/in2 0.03fF
C1668 addersubtractor_0/fulladder_1/XOR_0/NAND_1/w_32_0# addersubtractor_0/fulladder_1/XOR_0/NAND_3/in1 0.03fF
C1669 S0 A2 0.18fF
C1670 addersubtractor_0/fulladder_0/XOR_1/NAND_2/a_6_n14# gnd 0.59fF
C1671 vdd addersubtractor_0/fulladder_0/XOR_1/NAND_2/w_32_0# 0.05fF
C1672 XOR_0/NAND_2/a_6_n14# XOR_0/NAND_3/in2 0.12fF
C1673 vdd enableblock_2/enable1_0/AND_0/NAND_0/w_32_0# 0.05fF
C1674 vdd addersubtractor_0/fulladder_1/AND_0/not_0/in 0.29fF
C1675 addersubtractor_0/fulladder_0/XOR_1/NAND_1/w_0_0# S0 0.06fF
C1676 addersubtractor_0/fulladder_0/AND_1/not_0/w_0_0# addersubtractor_0/fulladder_0/AND_1/not_0/in 0.06fF
C1677 comparator_0/fiveinputAND_0/fiveinputNAND_0/w_0_0# comparator_0/fiveinputAND_0/not_0/in 0.03fF
C1678 vdd comparator_0/not_2/w_0_0# 0.05fF
C1679 enableblock_0/enable1_1/AND_1/not_0/w_0_0# enableblock_0/enable1_1/AND_1/not_0/in 0.06fF
C1680 vdd comparator_0/B0 0.17fF
C1681 vdd enableblock_1/enable1_0/AND_2/NAND_0/w_0_0# 0.05fF
C1682 addersubtractor_0/fulladder_0/XOR_0/NAND_2/a_6_n14# gnd 0.59fF
C1683 addersubtractor_0/fulladder_0/XOR_0/NAND_2/w_32_0# vdd 0.05fF
C1684 addersubtractor_0/fulladder_0/XOR_0/NAND_0/w_0_0# vdd 0.05fF
C1685 addersubtractor_0/fulladder_1/XOR_0/NAND_2/w_0_0# addersubtractor_0/fulladder_1/XOR_0/NAND_3/in2 0.03fF
C1686 enableblock_0/A_out1 gnd 1.72fF
C1687 addersubtractor_0/fulladder_2/XOR_0/NAND_2/in1 gnd 0.15fF
C1688 vdd addersubtractor_0/fulladder_2/AND_0/NAND_0/w_0_0# 0.05fF
C1689 comparator_0/fourinputOR_0/not_0/in comparator_0/fourinputOR_0/in2 0.11fF
C1690 addersubtractor_0/XOR_1/NAND_2/w_0_0# addersubtractor_0/XOR_1/NAND_3/in2 0.03fF
C1691 addersubtractor_0/fulladder_1/OR_0/NOT_0/in addersubtractor_0/fulladder_1/C 0.02fF
C1692 gnd AND_2/in1 0.16fF
C1693 AND_2/in2 enableblock_1/enable1_1/AND_3/NAND_0/w_0_0# 0.06fF
C1694 vdd addersubtractor_0/fulladder_3/AND_1/NAND_0/w_0_0# 0.05fF
C1695 vdd OR_0/NOR_0/w_0_0# 0.05fF
C1696 andblock_0/AND_1/NAND_0/a_6_n14# andblock_0/AND_1/not_0/in 0.12fF
C1697 vdd comparator_0/XNOR_0/not_0/w_0_0# 0.05fF
C1698 addersubtractor_0/fulladder_3/AND_0/not_0/in gnd 0.04fF
C1699 comparator_0/not_2/out comparator_0/B1 0.02fF
C1700 andblock_0/B2 enableblock_2/enable1_0/AND_3/not_0/in 0.02fF
C1701 OR_0/out enableblock_0/enable1_0/AND_2/NAND_0/w_32_0# 0.06fF
C1702 vdd addersubtractor_0/fulladder_1/OR_0/NOR_0/a_13_6# 0.21fF
C1703 addersubtractor_0/fulladder_1/OR_0/in1 gnd 0.30fF
C1704 gnd comparator_0/threeinputAND_0/threeinputNAND_0/a_45_n14# 0.04fF
C1705 vdd greater 0.39fF
C1706 addersubtractor_0/fulladder_3/AND_0/not_0/w_0_0# addersubtractor_0/fulladder_3/AND_0/not_0/in 0.06fF
C1707 vdd addersubtractor_0/XOR_1/out 0.32fF
C1708 gnd equal 0.08fF
C1709 vdd addersubtractor_0/fulladder_2/XOR_0/NAND_0/w_32_0# 0.05fF
C1710 vdd comparator_0/fourinputOR_0/in3 0.18fF
C1711 comparator_0/not_2/w_0_0# comparator_0/not_2/out 0.03fF
C1712 twotofourdecoder_0/AND_0/NAND_0/w_32_0# twotofourdecoder_0/AND_0/not_0/in 0.03fF
C1713 B2 B3 0.19fF
C1714 comparator_0/XNOR_1/XOR_0/NAND_0/w_0_0# comparator_0/XNOR_1/XOR_0/NAND_2/in1 0.03fF
C1715 enableblock_0/B_out1 enableblock_0/enable1_1/AND_2/not_0/w_0_0# 0.03fF
C1716 vdd addersubtractor_0/fulladder_2/XOR_1/NAND_0/w_32_0# 0.05fF
C1717 equal AND_2/not_0/w_0_0# 0.03fF
C1718 comparator_0/XNOR_2/out comparator_0/XNOR_2/not_0/in 0.02fF
C1719 comparator_0/AND_0/out comparator_0/AND_0/not_0/in 0.02fF
C1720 vdd comparator_0/fourinputOR_0/fourinputNOR_0/w_0_0# 0.05fF
C1721 vdd enableblock_0/B_out0 0.11fF
C1722 vdd addersubtractor_0/XOR_0/NAND_2/in1 0.25fF
C1723 vdd enableblock_1/enable1_0/AND_0/NAND_0/w_32_0# 0.05fF
C1724 S0 A3 0.20fF
C1725 gnd enableblock_1/enable1_1/AND_2/not_0/in 0.04fF
C1726 addersubtractor_0/fulladder_2/C addersubtractor_0/fulladder_3/XOR_1/NAND_1/w_0_0# 0.06fF
C1727 gnd addersubtractor_0/XOR_3/out 0.56fF
C1728 addersubtractor_0/fulladder_2/AND_1/NAND_0/w_32_0# addersubtractor_0/fulladder_2/AND_1/not_0/in 0.03fF
C1729 gnd comparator_0/A3 1.24fF
C1730 enableblock_1/enable1_0/AND_1/not_0/in comparator_0/B3 0.02fF
C1731 vdd addersubtractor_0/XOR_0/NAND_0/w_32_0# 0.05fF
C1732 AND_2/in2 lesser 0.06fF
C1733 AND_2/in2 A2 0.06fF
C1734 twotofourdecoder_0/AND_2/NAND_0/a_6_n14# twotofourdecoder_0/AND_2/not_0/in 0.12fF
C1735 vdd addersubtractor_0/fulladder_3/OR_0/NOT_0/w_0_0# 0.05fF
C1736 gnd comparator_0/A1 1.67fF
C1737 addersubtractor_0/fulladder_1/AND_0/not_0/in addersubtractor_0/fulladder_1/AND_0/NAND_0/a_6_n14# 0.12fF
C1738 vdd comparator_0/XNOR_0/XOR_0/NAND_0/w_0_0# 0.05fF
C1739 vdd andblock_0/B3 0.26fF
C1740 addersubtractor_0/XOR_2/NAND_0/w_0_0# enableblock_0/B_out2 0.06fF
C1741 gnd comparator_0/A0 1.10fF
C1742 vdd addersubtractor_0/XOR_3/NAND_0/w_0_0# 0.05fF
C1743 comparator_0/fourinputOR_0/in4 AND_2/in1 1.13fF
C1744 vdd comparator_0/XNOR_2/XOR_0/NAND_0/w_0_0# 0.05fF
C1745 andblock_0/AND_2/not_0/in andblock_0/AND_2/not_0/w_0_0# 0.06fF
C1746 OR_0/in2 OR_0/in1 0.06fF
C1747 addersubtractor_0/fulladder_1/AND_0/NAND_0/a_6_n14# addersubtractor_0/XOR_1/out 0.07fF
C1748 gnd comparator_0/AND_0/NAND_0/a_6_n14# 0.57fF
C1749 gnd enableblock_0/enable1_1/AND_1/NAND_0/a_6_n14# 0.57fF
C1750 vdd OR_0/out 0.13fF
C1751 vdd comparator_0/XNOR_3/XOR_0/NAND_0/w_0_0# 0.05fF
C1752 vdd addersubtractor_0/XOR_1/NAND_3/in2 0.25fF
C1753 OR_0/out B3 0.10fF
C1754 addersubtractor_0/fulladder_1/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_1/XOR_0/NAND_2/w_0_0# 0.06fF
C1755 vdd comparator_0/NOR_0/a_13_6# 0.21fF
C1756 vdd twotofourdecoder_0/AND_2/NAND_0/w_32_0# 0.05fF
C1757 gnd enableblock_0/enable1_0/AND_3/not_0/in 0.04fF
C1758 enableblock_1/enable1_0/AND_3/NAND_0/w_0_0# enableblock_1/enable1_0/AND_3/not_0/in 0.03fF
C1759 addersubtractor_0/XOR_3/NAND_1/w_0_0# enableblock_0/B_out0 0.06fF
C1760 addersubtractor_0/fulladder_0/OR_0/NOT_0/in gnd 0.60fF
C1761 enableblock_2/enable1_0/AND_2/not_0/w_0_0# enableblock_2/enable1_0/AND_2/not_0/in 0.06fF
C1762 comparator_0/fourinputOR_0/not_0/in greater 0.02fF
C1763 addersubtractor_0/fulladder_1/XOR_1/NAND_3/in1 gnd 0.11fF
C1764 enableblock_0/A_out1 addersubtractor_0/fulladder_1/XOR_0/NAND_0/w_0_0# 0.06fF
C1765 vdd addersubtractor_0/fulladder_1/XOR_1/NAND_1/w_0_0# 0.05fF
C1766 enableblock_2/En twotofourdecoder_0/AND_0/not_0/in 0.11fF
C1767 vdd enableblock_1/enable1_0/AND_2/not_0/in 0.29fF
C1768 addersubtractor_0/XOR_3/NAND_1/a_6_n14# addersubtractor_0/XOR_3/NAND_3/in1 0.12fF
C1769 B0 enableblock_2/En 0.06fF
C1770 comparator_0/B3 comparator_0/XNOR_0/XOR_0/NAND_2/w_32_0# 0.06fF
C1771 comparator_0/fourinputOR_0/not_0/in comparator_0/fourinputOR_0/in3 0.15fF
C1772 vdd addersubtractor_0/XOR_2/NAND_1/w_0_0# 0.05fF
C1773 addersubtractor_0/fulladder_1/XOR_0/NAND_3/in1 gnd 0.11fF
C1774 gnd andblock_0/AND_2/not_0/in 0.04fF
C1775 vdd addersubtractor_0/fulladder_1/XOR_0/NAND_1/w_0_0# 0.05fF
C1776 gnd enableblock_0/enable1_1/AND_2/NAND_0/a_6_n14# 0.57fF
C1777 S0 addersubtractor_0/XOR_2/NAND_0/w_32_0# 0.06fF
C1778 addersubtractor_0/fulladder_0/C addersubtractor_0/fulladder_1/XOR_1/in2 0.06fF
C1779 vdd enableblock_0/enable1_1/AND_1/not_0/w_0_0# 0.05fF
C1780 addersubtractor_0/fulladder_3/AND_0/not_0/in addersubtractor_0/fulladder_3/AND_0/NAND_0/w_0_0# 0.03fF
C1781 comparator_0/fourinputAND_0/not_0/w_0_0# comparator_0/fourinputOR_0/in3 0.03fF
C1782 enableblock_0/enable1_1/AND_2/NAND_0/w_32_0# enableblock_0/enable1_1/AND_2/not_0/in 0.03fF
C1783 gnd addersubtractor_0/fulladder_2/XOR_1/NAND_1/a_6_n14# 0.57fF
C1784 vdd addersubtractor_0/fulladder_2/XOR_1/NAND_1/w_32_0# 0.05fF
C1785 gnd comparator_0/AND_0/out 0.54fF
C1786 vdd enableblock_2/enable1_1/AND_3/NAND_0/w_0_0# 0.05fF
C1787 enableblock_0/A_out2 enableblock_0/enable1_0/AND_1/not_0/in 0.02fF
C1788 addersubtractor_0/fulladder_2/XOR_0/NAND_1/a_6_n14# gnd 0.57fF
C1789 vdd addersubtractor_0/fulladder_2/XOR_0/NAND_1/w_32_0# 0.05fF
C1790 addersubtractor_0/fulladder_1/OR_0/NOT_0/in addersubtractor_0/fulladder_1/OR_0/NOR_0/w_32_0# 0.03fF
C1791 comparator_0/B1 comparator_0/XNOR_2/XOR_0/NAND_2/w_32_0# 0.06fF
C1792 enableblock_0/enable1_1/AND_3/not_0/w_0_0# enableblock_0/B_out0 0.03fF
C1793 addersubtractor_0/XOR_2/out addersubtractor_0/fulladder_2/XOR_0/NAND_2/w_32_0# 0.06fF
C1794 gnd S0 1.94fF
C1795 vdd andblock_0/AND_0/NAND_0/w_32_0# 0.05fF
C1796 addersubtractor_0/fulladder_3/XOR_0/NAND_2/in1 addersubtractor_0/fulladder_3/XOR_0/NAND_0/a_6_n14# 0.12fF
C1797 addersubtractor_0/fulladder_3/AND_0/NAND_0/w_0_0# addersubtractor_0/XOR_3/out 0.06fF
C1798 addersubtractor_0/fulladder_3/AND_0/NAND_0/w_32_0# enableblock_0/B_out1 0.06fF
C1799 twotofourdecoder_0/AND_1/NAND_0/w_0_0# twotofourdecoder_0/AND_1/not_0/in 0.03fF
C1800 vdd addersubtractor_0/XOR_3/NAND_3/w_0_0# 0.05fF
C1801 comparator_0/B0 comparator_0/XNOR_3/XOR_0/NAND_2/w_32_0# 0.06fF
C1802 addersubtractor_0/fulladder_3/XOR_1/NAND_3/in1 addersubtractor_0/fulladder_3/XOR_1/NAND_3/w_0_0# 0.06fF
C1803 enableblock_1/enable1_1/AND_0/NAND_0/w_0_0# enableblock_1/enable1_1/AND_0/not_0/in 0.03fF
C1804 addersubtractor_0/fulladder_3/XOR_0/NAND_0/w_32_0# addersubtractor_0/XOR_3/out 0.06fF
C1805 addersubtractor_0/fulladder_0/XOR_1/NAND_0/w_0_0# S0 0.06fF
C1806 enableblock_1/enable1_1/AND_2/not_0/w_0_0# enableblock_1/enable1_1/AND_2/not_0/in 0.06fF
C1807 andblock_0/A0 andblock_0/AND_3/NAND_0/w_0_0# 0.06fF
C1808 addersubtractor_0/XOR_3/NAND_2/w_32_0# addersubtractor_0/XOR_3/NAND_3/in2 0.03fF
C1809 addersubtractor_0/XOR_1/out addersubtractor_0/XOR_1/NAND_3/w_0_0# 0.03fF
C1810 addersubtractor_0/fulladder_3/XOR_0/NAND_3/in1 addersubtractor_0/fulladder_3/XOR_0/NAND_3/w_0_0# 0.06fF
C1811 gnd enableblock_2/enable1_0/AND_3/NAND_0/a_6_n14# 0.57fF
C1812 vdd enableblock_2/enable1_0/AND_2/not_0/w_0_0# 0.05fF
C1813 addersubtractor_0/fulladder_3/AND_1/not_0/in addersubtractor_0/fulladder_3/OR_0/in1 0.02fF
C1814 A1 S1 0.06fF
C1815 gnd OR_0/NOT_0/in 0.60fF
C1816 enableblock_2/enable1_0/AND_1/NAND_0/a_6_n14# enableblock_2/enable1_0/AND_1/not_0/in 0.12fF
C1817 gnd enableblock_0/A_out2 0.92fF
C1818 enableblock_2/enable1_0/AND_0/not_0/in andblock_0/A3 0.02fF
C1819 gnd addersubtractor_0/XOR_1/NAND_2/a_6_n14# 0.59fF
C1820 vdd addersubtractor_0/XOR_1/NAND_2/w_32_0# 0.05fF
C1821 twotofourdecoder_0/AND_3/not_0/w_0_0# OR_0/in1 0.03fF
C1822 comparator_0/A3 comparator_0/XNOR_0/XOR_0/NAND_1/w_0_0# 0.06fF
C1823 comparator_0/XNOR_1/XOR_0/NAND_3/in1 comparator_0/XNOR_1/XOR_0/NAND_3/w_0_0# 0.06fF
C1824 addersubtractor_0/fulladder_3/OR_0/NOR_0/w_0_0# addersubtractor_0/fulladder_3/OR_0/in1 0.06fF
C1825 enableblock_1/enable1_1/AND_2/not_0/w_0_0# comparator_0/A0 0.03fF
C1826 enableblock_2/enable1_0/AND_1/not_0/w_0_0# andblock_0/B3 0.03fF
C1827 OR_0/NOR_0/a_13_6# Gnd 0.02fF
C1828 OR_0/NOR_0/w_32_0# Gnd 0.40fF
C1829 OR_0/NOR_0/w_0_0# Gnd 0.40fF
C1830 OR_0/NOT_0/in Gnd 0.77fF
C1831 OR_0/NOT_0/w_0_0# Gnd 0.40fF
C1832 XOR_0/NAND_3/a_6_n14# Gnd 0.14fF
C1833 Carry Gnd 0.53fF
C1834 XOR_0/NAND_3/in2 Gnd 0.76fF
C1835 XOR_0/NAND_3/w_32_0# Gnd 0.40fF
C1836 XOR_0/NAND_3/w_0_0# Gnd 0.40fF
C1837 XOR_0/NAND_2/a_6_n14# Gnd 0.14fF
C1838 XOR_0/NAND_2/w_32_0# Gnd 0.40fF
C1839 XOR_0/NAND_2/w_0_0# Gnd 0.40fF
C1840 XOR_0/NAND_1/a_6_n14# Gnd 0.14fF
C1841 XOR_0/NAND_3/in1 Gnd 0.78fF
C1842 XOR_0/NAND_1/w_32_0# Gnd 0.40fF
C1843 XOR_0/NAND_1/w_0_0# Gnd 0.40fF
C1844 XOR_0/NAND_0/a_6_n14# Gnd 0.14fF
C1845 XOR_0/NAND_2/in1 Gnd 0.97fF
C1846 XOR_0/in1 Gnd 1.72fF
C1847 XOR_0/NAND_0/w_32_0# Gnd 0.40fF
C1848 XOR_0/NAND_0/w_0_0# Gnd 0.40fF
C1849 andblock_0/AND_3/not_0/in Gnd 0.76fF
C1850 and0 Gnd 0.19fF
C1851 andblock_0/AND_3/not_0/w_0_0# Gnd 0.40fF
C1852 andblock_0/AND_3/NAND_0/a_6_n14# Gnd 0.14fF
C1853 andblock_0/AND_3/NAND_0/w_32_0# Gnd 0.40fF
C1854 andblock_0/AND_3/NAND_0/w_0_0# Gnd 0.40fF
C1855 andblock_0/AND_2/not_0/in Gnd 0.76fF
C1856 and1 Gnd 0.20fF
C1857 andblock_0/AND_2/not_0/w_0_0# Gnd 0.40fF
C1858 andblock_0/AND_2/NAND_0/a_6_n14# Gnd 0.14fF
C1859 andblock_0/AND_2/NAND_0/w_32_0# Gnd 0.40fF
C1860 andblock_0/AND_2/NAND_0/w_0_0# Gnd 0.40fF
C1861 andblock_0/AND_1/not_0/in Gnd 0.76fF
C1862 and2 Gnd 0.20fF
C1863 andblock_0/AND_1/not_0/w_0_0# Gnd 0.40fF
C1864 andblock_0/AND_1/NAND_0/a_6_n14# Gnd 0.14fF
C1865 andblock_0/AND_1/NAND_0/w_32_0# Gnd 0.40fF
C1866 andblock_0/AND_1/NAND_0/w_0_0# Gnd 0.40fF
C1867 andblock_0/AND_0/not_0/in Gnd 0.76fF
C1868 and3 Gnd 0.20fF
C1869 andblock_0/AND_0/not_0/w_0_0# Gnd 0.40fF
C1870 andblock_0/AND_0/NAND_0/a_6_n14# Gnd 0.14fF
C1871 andblock_0/AND_0/NAND_0/w_32_0# Gnd 0.40fF
C1872 andblock_0/AND_0/NAND_0/w_0_0# Gnd 0.40fF
C1873 lesser Gnd 0.67fF
C1874 comparator_0/NOR_0/a_13_6# Gnd 0.02fF
C1875 comparator_0/NOR_0/w_32_0# Gnd 0.40fF
C1876 comparator_0/NOR_0/w_0_0# Gnd 0.40fF
C1877 comparator_0/XNOR_3/XOR_0/NAND_3/a_6_n14# Gnd 0.14fF
C1878 comparator_0/XNOR_3/not_0/in Gnd 0.76fF
C1879 comparator_0/XNOR_3/XOR_0/NAND_3/in2 Gnd 0.76fF
C1880 comparator_0/XNOR_3/XOR_0/NAND_3/w_32_0# Gnd 0.40fF
C1881 comparator_0/XNOR_3/XOR_0/NAND_3/w_0_0# Gnd 0.40fF
C1882 comparator_0/XNOR_3/XOR_0/NAND_2/a_6_n14# Gnd 0.14fF
C1883 comparator_0/XNOR_3/XOR_0/NAND_2/w_32_0# Gnd 0.40fF
C1884 comparator_0/XNOR_3/XOR_0/NAND_2/w_0_0# Gnd 0.40fF
C1885 comparator_0/XNOR_3/XOR_0/NAND_1/a_6_n14# Gnd 0.14fF
C1886 comparator_0/XNOR_3/XOR_0/NAND_3/in1 Gnd 0.78fF
C1887 comparator_0/XNOR_3/XOR_0/NAND_1/w_32_0# Gnd 0.40fF
C1888 comparator_0/XNOR_3/XOR_0/NAND_1/w_0_0# Gnd 0.40fF
C1889 comparator_0/XNOR_3/XOR_0/NAND_0/a_6_n14# Gnd 0.14fF
C1890 comparator_0/XNOR_3/XOR_0/NAND_2/in1 Gnd 0.97fF
C1891 comparator_0/B0 Gnd 1.82fF
C1892 comparator_0/A0 Gnd 3.08fF
C1893 comparator_0/XNOR_3/XOR_0/NAND_0/w_32_0# Gnd 0.40fF
C1894 comparator_0/XNOR_3/XOR_0/NAND_0/w_0_0# Gnd 0.40fF
C1895 comparator_0/XNOR_3/not_0/w_0_0# Gnd 0.40fF
C1896 comparator_0/XNOR_2/XOR_0/NAND_3/a_6_n14# Gnd 0.14fF
C1897 comparator_0/XNOR_2/not_0/in Gnd 0.76fF
C1898 comparator_0/XNOR_2/XOR_0/NAND_3/in2 Gnd 0.76fF
C1899 comparator_0/XNOR_2/XOR_0/NAND_3/w_32_0# Gnd 0.40fF
C1900 comparator_0/XNOR_2/XOR_0/NAND_3/w_0_0# Gnd 0.40fF
C1901 comparator_0/XNOR_2/XOR_0/NAND_2/a_6_n14# Gnd 0.14fF
C1902 comparator_0/XNOR_2/XOR_0/NAND_2/w_32_0# Gnd 0.40fF
C1903 comparator_0/XNOR_2/XOR_0/NAND_2/w_0_0# Gnd 0.40fF
C1904 comparator_0/XNOR_2/XOR_0/NAND_1/a_6_n14# Gnd 0.14fF
C1905 comparator_0/XNOR_2/XOR_0/NAND_3/in1 Gnd 0.78fF
C1906 comparator_0/XNOR_2/XOR_0/NAND_1/w_32_0# Gnd 0.40fF
C1907 comparator_0/XNOR_2/XOR_0/NAND_1/w_0_0# Gnd 0.40fF
C1908 comparator_0/XNOR_2/XOR_0/NAND_0/a_6_n14# Gnd 0.14fF
C1909 comparator_0/XNOR_2/XOR_0/NAND_2/in1 Gnd 0.97fF
C1910 comparator_0/B1 Gnd 1.62fF
C1911 comparator_0/A1 Gnd 2.60fF
C1912 comparator_0/XNOR_2/XOR_0/NAND_0/w_32_0# Gnd 0.40fF
C1913 comparator_0/XNOR_2/XOR_0/NAND_0/w_0_0# Gnd 0.40fF
C1914 comparator_0/XNOR_2/not_0/w_0_0# Gnd 0.40fF
C1915 comparator_0/XNOR_0/XOR_0/NAND_3/a_6_n14# Gnd 0.14fF
C1916 comparator_0/XNOR_0/not_0/in Gnd 0.76fF
C1917 comparator_0/XNOR_0/XOR_0/NAND_3/in2 Gnd 0.76fF
C1918 comparator_0/XNOR_0/XOR_0/NAND_3/w_32_0# Gnd 0.40fF
C1919 comparator_0/XNOR_0/XOR_0/NAND_3/w_0_0# Gnd 0.40fF
C1920 comparator_0/XNOR_0/XOR_0/NAND_2/a_6_n14# Gnd 0.14fF
C1921 comparator_0/XNOR_0/XOR_0/NAND_2/w_32_0# Gnd 0.40fF
C1922 comparator_0/XNOR_0/XOR_0/NAND_2/w_0_0# Gnd 0.40fF
C1923 comparator_0/XNOR_0/XOR_0/NAND_1/a_6_n14# Gnd 0.14fF
C1924 comparator_0/XNOR_0/XOR_0/NAND_3/in1 Gnd 0.78fF
C1925 comparator_0/XNOR_0/XOR_0/NAND_1/w_32_0# Gnd 0.40fF
C1926 comparator_0/XNOR_0/XOR_0/NAND_1/w_0_0# Gnd 0.40fF
C1927 comparator_0/XNOR_0/XOR_0/NAND_0/a_6_n14# Gnd 0.14fF
C1928 comparator_0/XNOR_0/XOR_0/NAND_2/in1 Gnd 0.97fF
C1929 comparator_0/B3 Gnd 0.01fF
C1930 comparator_0/A3 Gnd 1.29fF
C1931 comparator_0/XNOR_0/XOR_0/NAND_0/w_32_0# Gnd 0.40fF
C1932 comparator_0/XNOR_0/XOR_0/NAND_0/w_0_0# Gnd 0.40fF
C1933 comparator_0/XNOR_0/not_0/w_0_0# Gnd 0.40fF
C1934 comparator_0/XNOR_1/XOR_0/NAND_3/a_6_n14# Gnd 0.14fF
C1935 comparator_0/XNOR_1/not_0/in Gnd 0.76fF
C1936 comparator_0/XNOR_1/XOR_0/NAND_3/in2 Gnd 0.76fF
C1937 comparator_0/XNOR_1/XOR_0/NAND_3/w_32_0# Gnd 0.40fF
C1938 comparator_0/XNOR_1/XOR_0/NAND_3/w_0_0# Gnd 0.40fF
C1939 comparator_0/XNOR_1/XOR_0/NAND_2/a_6_n14# Gnd 0.14fF
C1940 comparator_0/XNOR_1/XOR_0/NAND_2/w_32_0# Gnd 0.40fF
C1941 comparator_0/XNOR_1/XOR_0/NAND_2/w_0_0# Gnd 0.40fF
C1942 comparator_0/XNOR_1/XOR_0/NAND_1/a_6_n14# Gnd 0.14fF
C1943 comparator_0/XNOR_1/XOR_0/NAND_3/in1 Gnd 0.78fF
C1944 comparator_0/XNOR_1/XOR_0/NAND_1/w_32_0# Gnd 0.40fF
C1945 comparator_0/XNOR_1/XOR_0/NAND_1/w_0_0# Gnd 0.40fF
C1946 comparator_0/XNOR_1/XOR_0/NAND_0/a_6_n14# Gnd 0.14fF
C1947 comparator_0/XNOR_1/XOR_0/NAND_2/in1 Gnd 0.97fF
C1948 comparator_0/B2 Gnd 2.68fF
C1949 comparator_0/A2 Gnd 2.23fF
C1950 comparator_0/XNOR_1/XOR_0/NAND_0/w_32_0# Gnd 0.40fF
C1951 comparator_0/XNOR_1/XOR_0/NAND_0/w_0_0# Gnd 0.40fF
C1952 comparator_0/XNOR_1/not_0/w_0_0# Gnd 0.40fF
C1953 comparator_0/fiveinputAND_0/fiveinputNAND_0/a_113_n14# Gnd 0.08fF
C1954 comparator_0/fiveinputAND_0/fiveinputNAND_0/a_76_n14# Gnd 0.05fF
C1955 comparator_0/fiveinputAND_0/fiveinputNAND_0/a_45_n14# Gnd 0.07fF
C1956 comparator_0/fiveinputAND_0/fiveinputNAND_0/a_6_n14# Gnd 0.14fF
C1957 comparator_0/XNOR_2/out Gnd 1.52fF
C1958 comparator_0/not_3/out Gnd 1.44fF
C1959 comparator_0/fiveinputAND_0/fiveinputNAND_0/w_133_0# Gnd 0.43fF
C1960 comparator_0/fiveinputAND_0/fiveinputNAND_0/w_63_0# Gnd 0.43fF
C1961 comparator_0/fiveinputAND_0/fiveinputNAND_0/w_32_0# Gnd 0.43fF
C1962 comparator_0/fiveinputAND_0/fiveinputNAND_0/w_0_0# Gnd 0.43fF
C1963 comparator_0/fiveinputAND_0/not_0/in Gnd 1.48fF
C1964 comparator_0/fiveinputAND_0/not_0/w_0_0# Gnd 0.40fF
C1965 comparator_0/fourinputOR_0/in2 Gnd 1.03fF
C1966 comparator_0/threeinputAND_0/not_0/in Gnd 0.76fF
C1967 comparator_0/threeinputAND_0/not_0/w_0_0# Gnd 0.40fF
C1968 comparator_0/threeinputAND_0/threeinputNAND_0/a_45_n14# Gnd 0.07fF
C1969 comparator_0/threeinputAND_0/threeinputNAND_0/a_6_n14# Gnd 0.14fF
C1970 comparator_0/XNOR_0/out Gnd 0.53fF
C1971 comparator_0/not_1/out Gnd 0.29fF
C1972 comparator_0/threeinputAND_0/threeinputNAND_0/w_63_0# Gnd 0.39fF
C1973 comparator_0/threeinputAND_0/threeinputNAND_0/w_32_0# Gnd 0.40fF
C1974 comparator_0/threeinputAND_0/threeinputNAND_0/w_0_0# Gnd 0.40fF
C1975 comparator_0/fourinputAND_1/fourinputNAND_0/a_76_n14# Gnd 0.05fF
C1976 comparator_0/fourinputAND_1/fourinputNAND_0/a_45_n14# Gnd 0.07fF
C1977 comparator_0/fourinputAND_1/fourinputNAND_0/a_6_n14# Gnd 0.14fF
C1978 comparator_0/fourinputAND_1/not_0/in Gnd 1.84fF
C1979 comparator_0/XNOR_3/out Gnd 0.61fF
C1980 comparator_0/fourinputAND_1/fourinputNAND_0/w_100_0# Gnd 0.40fF
C1981 comparator_0/fourinputAND_1/fourinputNAND_0/w_63_0# Gnd 0.40fF
C1982 comparator_0/fourinputAND_1/fourinputNAND_0/w_32_0# Gnd 0.40fF
C1983 comparator_0/fourinputAND_1/fourinputNAND_0/w_0_0# Gnd 0.40fF
C1984 comparator_0/fourinputAND_1/not_0/w_0_0# Gnd 0.40fF
C1985 comparator_0/fourinputAND_0/fourinputNAND_0/a_76_n14# Gnd 0.05fF
C1986 comparator_0/fourinputAND_0/fourinputNAND_0/a_45_n14# Gnd 0.07fF
C1987 comparator_0/fourinputAND_0/fourinputNAND_0/a_6_n14# Gnd 0.14fF
C1988 comparator_0/fourinputAND_0/not_0/in Gnd 1.84fF
C1989 comparator_0/not_2/out Gnd 0.30fF
C1990 comparator_0/fourinputAND_0/fourinputNAND_0/w_100_0# Gnd 0.40fF
C1991 comparator_0/fourinputAND_0/fourinputNAND_0/w_63_0# Gnd 0.40fF
C1992 comparator_0/fourinputAND_0/fourinputNAND_0/w_32_0# Gnd 0.40fF
C1993 comparator_0/fourinputAND_0/fourinputNAND_0/w_0_0# Gnd 0.40fF
C1994 comparator_0/fourinputOR_0/in3 Gnd 1.03fF
C1995 comparator_0/fourinputAND_0/not_0/w_0_0# Gnd 0.40fF
C1996 comparator_0/not_3/w_0_0# Gnd 0.40fF
C1997 comparator_0/not_2/w_0_0# Gnd 0.40fF
C1998 comparator_0/not_1/w_0_0# Gnd 0.40fF
C1999 comparator_0/not_0/w_0_0# Gnd 0.40fF
C2000 comparator_0/AND_0/not_0/in Gnd 0.76fF
C2001 comparator_0/AND_0/out Gnd 1.01fF
C2002 comparator_0/AND_0/not_0/w_0_0# Gnd 0.40fF
C2003 comparator_0/AND_0/NAND_0/a_6_n14# Gnd 0.14fF
C2004 comparator_0/not_0/out Gnd 0.28fF
C2005 comparator_0/AND_0/NAND_0/w_32_0# Gnd 0.40fF
C2006 comparator_0/AND_0/NAND_0/w_0_0# Gnd 0.40fF
C2007 greater Gnd 1.58fF
C2008 comparator_0/fourinputOR_0/not_0/in Gnd 1.09fF
C2009 comparator_0/fourinputOR_0/not_0/w_0_0# Gnd 0.40fF
C2010 comparator_0/fourinputOR_0/fourinputNOR_0/a_77_6# Gnd 0.02fF
C2011 comparator_0/fourinputOR_0/fourinputNOR_0/a_45_6# Gnd 0.02fF
C2012 comparator_0/fourinputOR_0/fourinputNOR_0/a_13_6# Gnd 0.02fF
C2013 comparator_0/fourinputOR_0/in4 Gnd 0.13fF
C2014 comparator_0/fourinputOR_0/fourinputNOR_0/w_97_0# Gnd 0.03fF
C2015 comparator_0/fourinputOR_0/fourinputNOR_0/w_64_0# Gnd 0.40fF
C2016 comparator_0/fourinputOR_0/fourinputNOR_0/w_32_0# Gnd 0.40fF
C2017 comparator_0/fourinputOR_0/fourinputNOR_0/w_0_0# Gnd 0.40fF
C2018 twotofourdecoder_0/not_1/w_0_0# Gnd 0.40fF
C2019 twotofourdecoder_0/not_0/w_0_0# Gnd 0.40fF
C2020 twotofourdecoder_0/AND_3/not_0/in Gnd 0.76fF
C2021 twotofourdecoder_0/AND_3/not_0/w_0_0# Gnd 0.40fF
C2022 twotofourdecoder_0/AND_3/NAND_0/a_6_n14# Gnd 0.14fF
C2023 twotofourdecoder_0/not_1/out Gnd 1.39fF
C2024 twotofourdecoder_0/AND_3/NAND_0/w_32_0# Gnd 0.40fF
C2025 twotofourdecoder_0/AND_3/NAND_0/w_0_0# Gnd 0.40fF
C2026 twotofourdecoder_0/AND_2/not_0/in Gnd 0.76fF
C2027 OR_0/in2 Gnd 4.82fF
C2028 twotofourdecoder_0/AND_2/not_0/w_0_0# Gnd 0.40fF
C2029 twotofourdecoder_0/AND_2/NAND_0/a_6_n14# Gnd 0.14fF
C2030 twotofourdecoder_0/AND_2/NAND_0/w_32_0# Gnd 0.40fF
C2031 twotofourdecoder_0/AND_2/NAND_0/w_0_0# Gnd 0.40fF
C2032 twotofourdecoder_0/AND_1/not_0/in Gnd 0.76fF
C2033 twotofourdecoder_0/AND_1/not_0/w_0_0# Gnd 0.40fF
C2034 twotofourdecoder_0/AND_1/NAND_0/a_6_n14# Gnd 0.14fF
C2035 twotofourdecoder_0/not_0/out Gnd 1.67fF
C2036 twotofourdecoder_0/AND_1/NAND_0/w_32_0# Gnd 0.40fF
C2037 twotofourdecoder_0/AND_1/NAND_0/w_0_0# Gnd 0.40fF
C2038 twotofourdecoder_0/AND_0/not_0/in Gnd 0.76fF
C2039 twotofourdecoder_0/AND_0/not_0/w_0_0# Gnd 0.40fF
C2040 twotofourdecoder_0/AND_0/NAND_0/a_6_n14# Gnd 0.14fF
C2041 S1 Gnd 1.63fF
C2042 twotofourdecoder_0/AND_0/NAND_0/w_32_0# Gnd 0.40fF
C2043 twotofourdecoder_0/AND_0/NAND_0/w_0_0# Gnd 0.40fF
C2044 enableblock_2/enable1_1/AND_3/not_0/in Gnd 0.76fF
C2045 andblock_0/B0 Gnd 0.49fF
C2046 enableblock_2/enable1_1/AND_3/not_0/w_0_0# Gnd 0.40fF
C2047 enableblock_2/enable1_1/AND_3/NAND_0/a_6_n14# Gnd 0.14fF
C2048 enableblock_2/enable1_1/AND_3/NAND_0/w_32_0# Gnd 0.40fF
C2049 enableblock_2/enable1_1/AND_3/NAND_0/w_0_0# Gnd 0.40fF
C2050 enableblock_2/enable1_1/AND_2/not_0/in Gnd 0.76fF
C2051 andblock_0/A0 Gnd 0.33fF
C2052 enableblock_2/enable1_1/AND_2/not_0/w_0_0# Gnd 0.40fF
C2053 enableblock_2/enable1_1/AND_2/NAND_0/a_6_n14# Gnd 0.14fF
C2054 enableblock_2/enable1_1/AND_2/NAND_0/w_32_0# Gnd 0.40fF
C2055 enableblock_2/enable1_1/AND_2/NAND_0/w_0_0# Gnd 0.40fF
C2056 enableblock_2/enable1_1/AND_1/not_0/in Gnd 0.76fF
C2057 andblock_0/B1 Gnd 1.33fF
C2058 enableblock_2/enable1_1/AND_1/not_0/w_0_0# Gnd 0.40fF
C2059 enableblock_2/enable1_1/AND_1/NAND_0/a_6_n14# Gnd 0.14fF
C2060 enableblock_2/enable1_1/AND_1/NAND_0/w_32_0# Gnd 0.40fF
C2061 enableblock_2/enable1_1/AND_1/NAND_0/w_0_0# Gnd 0.40fF
C2062 enableblock_2/enable1_1/AND_0/not_0/in Gnd 0.76fF
C2063 andblock_0/A1 Gnd 0.86fF
C2064 enableblock_2/enable1_1/AND_0/not_0/w_0_0# Gnd 0.40fF
C2065 enableblock_2/enable1_1/AND_0/NAND_0/a_6_n14# Gnd 0.14fF
C2066 enableblock_2/enable1_1/AND_0/NAND_0/w_32_0# Gnd 0.40fF
C2067 enableblock_2/enable1_1/AND_0/NAND_0/w_0_0# Gnd 0.40fF
C2068 enableblock_2/enable1_0/AND_3/not_0/in Gnd 0.76fF
C2069 andblock_0/B2 Gnd 0.43fF
C2070 enableblock_2/enable1_0/AND_3/not_0/w_0_0# Gnd 0.40fF
C2071 enableblock_2/enable1_0/AND_3/NAND_0/a_6_n14# Gnd 0.14fF
C2072 enableblock_2/enable1_0/AND_3/NAND_0/w_32_0# Gnd 0.40fF
C2073 enableblock_2/enable1_0/AND_3/NAND_0/w_0_0# Gnd 0.40fF
C2074 enableblock_2/enable1_0/AND_2/not_0/in Gnd 0.76fF
C2075 andblock_0/A2 Gnd 0.78fF
C2076 enableblock_2/enable1_0/AND_2/not_0/w_0_0# Gnd 0.40fF
C2077 enableblock_2/enable1_0/AND_2/NAND_0/a_6_n14# Gnd 0.14fF
C2078 enableblock_2/enable1_0/AND_2/NAND_0/w_32_0# Gnd 0.40fF
C2079 enableblock_2/enable1_0/AND_2/NAND_0/w_0_0# Gnd 0.40fF
C2080 enableblock_2/enable1_0/AND_1/not_0/in Gnd 0.76fF
C2081 andblock_0/B3 Gnd 1.61fF
C2082 enableblock_2/enable1_0/AND_1/not_0/w_0_0# Gnd 0.40fF
C2083 enableblock_2/enable1_0/AND_1/NAND_0/a_6_n14# Gnd 0.14fF
C2084 enableblock_2/En Gnd 5.01fF
C2085 enableblock_2/enable1_0/AND_1/NAND_0/w_32_0# Gnd 0.40fF
C2086 enableblock_2/enable1_0/AND_1/NAND_0/w_0_0# Gnd 0.40fF
C2087 enableblock_2/enable1_0/AND_0/not_0/in Gnd 0.76fF
C2088 enableblock_2/enable1_0/AND_0/not_0/w_0_0# Gnd 0.40fF
C2089 enableblock_2/enable1_0/AND_0/NAND_0/a_6_n14# Gnd 0.14fF
C2090 enableblock_2/enable1_0/AND_0/NAND_0/w_32_0# Gnd 0.40fF
C2091 enableblock_2/enable1_0/AND_0/NAND_0/w_0_0# Gnd 0.40fF
C2092 enableblock_0/enable1_1/AND_3/not_0/in Gnd 0.76fF
C2093 enableblock_0/B_out0 Gnd 0.22fF
C2094 enableblock_0/enable1_1/AND_3/not_0/w_0_0# Gnd 0.40fF
C2095 enableblock_0/enable1_1/AND_3/NAND_0/a_6_n14# Gnd 0.14fF
C2096 B3 Gnd 40.94fF
C2097 enableblock_0/enable1_1/AND_3/NAND_0/w_32_0# Gnd 0.40fF
C2098 enableblock_0/enable1_1/AND_3/NAND_0/w_0_0# Gnd 0.40fF
C2099 enableblock_0/enable1_1/AND_2/not_0/in Gnd 0.76fF
C2100 enableblock_0/enable1_1/AND_2/not_0/w_0_0# Gnd 0.40fF
C2101 enableblock_0/enable1_1/AND_2/NAND_0/a_6_n14# Gnd 0.14fF
C2102 A3 Gnd 1.15fF
C2103 enableblock_0/enable1_1/AND_2/NAND_0/w_32_0# Gnd 0.40fF
C2104 enableblock_0/enable1_1/AND_2/NAND_0/w_0_0# Gnd 0.40fF
C2105 enableblock_0/enable1_1/AND_1/not_0/in Gnd 0.76fF
C2106 enableblock_0/B_out2 Gnd 1.70fF
C2107 enableblock_0/enable1_1/AND_1/not_0/w_0_0# Gnd 0.40fF
C2108 enableblock_0/enable1_1/AND_1/NAND_0/a_6_n14# Gnd 0.14fF
C2109 B2 Gnd 40.41fF
C2110 enableblock_0/enable1_1/AND_1/NAND_0/w_32_0# Gnd 0.40fF
C2111 enableblock_0/enable1_1/AND_1/NAND_0/w_0_0# Gnd 0.40fF
C2112 enableblock_0/enable1_1/AND_0/not_0/in Gnd 0.76fF
C2113 enableblock_0/enable1_1/AND_0/not_0/w_0_0# Gnd 0.40fF
C2114 enableblock_0/enable1_1/AND_0/NAND_0/a_6_n14# Gnd 0.14fF
C2115 A2 Gnd 39.38fF
C2116 enableblock_0/enable1_1/AND_0/NAND_0/w_32_0# Gnd 0.40fF
C2117 enableblock_0/enable1_1/AND_0/NAND_0/w_0_0# Gnd 0.40fF
C2118 enableblock_0/enable1_0/AND_3/not_0/in Gnd 0.76fF
C2119 enableblock_0/A_out0 Gnd 1.45fF
C2120 enableblock_0/enable1_0/AND_3/not_0/w_0_0# Gnd 0.40fF
C2121 enableblock_0/enable1_0/AND_3/NAND_0/a_6_n14# Gnd 0.14fF
C2122 B1 Gnd 40.05fF
C2123 enableblock_0/enable1_0/AND_3/NAND_0/w_32_0# Gnd 0.40fF
C2124 enableblock_0/enable1_0/AND_3/NAND_0/w_0_0# Gnd 0.40fF
C2125 enableblock_0/enable1_0/AND_2/not_0/in Gnd 0.76fF
C2126 enableblock_0/enable1_0/AND_2/not_0/w_0_0# Gnd 0.40fF
C2127 enableblock_0/enable1_0/AND_2/NAND_0/a_6_n14# Gnd 0.14fF
C2128 A1 Gnd 1.13fF
C2129 enableblock_0/enable1_0/AND_2/NAND_0/w_32_0# Gnd 0.40fF
C2130 enableblock_0/enable1_0/AND_2/NAND_0/w_0_0# Gnd 0.40fF
C2131 enableblock_0/enable1_0/AND_1/not_0/in Gnd 0.76fF
C2132 enableblock_0/A_out2 Gnd 1.63fF
C2133 enableblock_0/enable1_0/AND_1/not_0/w_0_0# Gnd 0.40fF
C2134 enableblock_0/enable1_0/AND_1/NAND_0/a_6_n14# Gnd 0.14fF
C2135 B0 Gnd 39.80fF
C2136 OR_0/out Gnd 5.23fF
C2137 enableblock_0/enable1_0/AND_1/NAND_0/w_32_0# Gnd 0.40fF
C2138 enableblock_0/enable1_0/AND_1/NAND_0/w_0_0# Gnd 0.40fF
C2139 enableblock_0/enable1_0/AND_0/not_0/in Gnd 0.76fF
C2140 enableblock_0/enable1_0/AND_0/not_0/w_0_0# Gnd 0.40fF
C2141 enableblock_0/enable1_0/AND_0/NAND_0/a_6_n14# Gnd 0.14fF
C2142 A0 Gnd 1.27fF
C2143 enableblock_0/enable1_0/AND_0/NAND_0/w_32_0# Gnd 0.40fF
C2144 enableblock_0/enable1_0/AND_0/NAND_0/w_0_0# Gnd 0.40fF
C2145 enableblock_1/enable1_1/AND_3/not_0/in Gnd 0.76fF
C2146 enableblock_1/enable1_1/AND_3/not_0/w_0_0# Gnd 0.40fF
C2147 enableblock_1/enable1_1/AND_3/NAND_0/a_6_n14# Gnd 0.14fF
C2148 enableblock_1/enable1_1/AND_3/NAND_0/w_32_0# Gnd 0.40fF
C2149 enableblock_1/enable1_1/AND_3/NAND_0/w_0_0# Gnd 0.40fF
C2150 enableblock_1/enable1_1/AND_2/not_0/in Gnd 0.76fF
C2151 enableblock_1/enable1_1/AND_2/not_0/w_0_0# Gnd 0.40fF
C2152 enableblock_1/enable1_1/AND_2/NAND_0/a_6_n14# Gnd 0.14fF
C2153 enableblock_1/enable1_1/AND_2/NAND_0/w_32_0# Gnd 0.40fF
C2154 enableblock_1/enable1_1/AND_2/NAND_0/w_0_0# Gnd 0.40fF
C2155 enableblock_1/enable1_1/AND_1/not_0/in Gnd 0.76fF
C2156 enableblock_1/enable1_1/AND_1/not_0/w_0_0# Gnd 0.40fF
C2157 enableblock_1/enable1_1/AND_1/NAND_0/a_6_n14# Gnd 0.14fF
C2158 enableblock_1/enable1_1/AND_1/NAND_0/w_32_0# Gnd 0.40fF
C2159 enableblock_1/enable1_1/AND_1/NAND_0/w_0_0# Gnd 0.40fF
C2160 enableblock_1/enable1_1/AND_0/not_0/in Gnd 0.76fF
C2161 enableblock_1/enable1_1/AND_0/not_0/w_0_0# Gnd 0.40fF
C2162 enableblock_1/enable1_1/AND_0/NAND_0/a_6_n14# Gnd 0.14fF
C2163 enableblock_1/enable1_1/AND_0/NAND_0/w_32_0# Gnd 0.40fF
C2164 enableblock_1/enable1_1/AND_0/NAND_0/w_0_0# Gnd 0.40fF
C2165 enableblock_1/enable1_0/AND_3/not_0/in Gnd 0.76fF
C2166 enableblock_1/enable1_0/AND_3/not_0/w_0_0# Gnd 0.40fF
C2167 enableblock_1/enable1_0/AND_3/NAND_0/a_6_n14# Gnd 0.14fF
C2168 enableblock_1/enable1_0/AND_3/NAND_0/w_32_0# Gnd 0.40fF
C2169 enableblock_1/enable1_0/AND_3/NAND_0/w_0_0# Gnd 0.40fF
C2170 enableblock_1/enable1_0/AND_2/not_0/in Gnd 0.76fF
C2171 enableblock_1/enable1_0/AND_2/not_0/w_0_0# Gnd 0.40fF
C2172 enableblock_1/enable1_0/AND_2/NAND_0/a_6_n14# Gnd 0.14fF
C2173 enableblock_1/enable1_0/AND_2/NAND_0/w_32_0# Gnd 0.40fF
C2174 enableblock_1/enable1_0/AND_2/NAND_0/w_0_0# Gnd 0.40fF
C2175 enableblock_1/enable1_0/AND_1/not_0/in Gnd 0.76fF
C2176 enableblock_1/enable1_0/AND_1/not_0/w_0_0# Gnd 0.40fF
C2177 enableblock_1/enable1_0/AND_1/NAND_0/a_6_n14# Gnd 0.14fF
C2178 AND_2/in2 Gnd 14.89fF
C2179 enableblock_1/enable1_0/AND_1/NAND_0/w_32_0# Gnd 0.40fF
C2180 enableblock_1/enable1_0/AND_1/NAND_0/w_0_0# Gnd 0.40fF
C2181 enableblock_1/enable1_0/AND_0/not_0/in Gnd 0.76fF
C2182 enableblock_1/enable1_0/AND_0/not_0/w_0_0# Gnd 0.40fF
C2183 enableblock_1/enable1_0/AND_0/NAND_0/a_6_n14# Gnd 0.14fF
C2184 enableblock_1/enable1_0/AND_0/NAND_0/w_32_0# Gnd 0.40fF
C2185 enableblock_1/enable1_0/AND_0/NAND_0/w_0_0# Gnd 0.40fF
C2186 AND_2/not_0/in Gnd 0.76fF
C2187 equal Gnd 0.17fF
C2188 AND_2/not_0/w_0_0# Gnd 0.40fF
C2189 AND_2/NAND_0/a_6_n14# Gnd 0.14fF
C2190 AND_2/NAND_0/w_32_0# Gnd 0.40fF
C2191 AND_2/NAND_0/w_0_0# Gnd 0.40fF
C2192 AND_0/not_0/in Gnd 0.76fF
C2193 AND_0/not_0/w_0_0# Gnd 0.40fF
C2194 AND_0/NAND_0/a_6_n14# Gnd 0.14fF
C2195 AND_0/NAND_0/w_32_0# Gnd 0.40fF
C2196 AND_0/NAND_0/w_0_0# Gnd 0.40fF
C2197 addersubtractor_0/XOR_3/NAND_3/a_6_n14# Gnd 0.14fF
C2198 addersubtractor_0/XOR_3/NAND_3/in2 Gnd 0.76fF
C2199 addersubtractor_0/XOR_3/NAND_3/w_32_0# Gnd 0.40fF
C2200 addersubtractor_0/XOR_3/NAND_3/w_0_0# Gnd 0.40fF
C2201 addersubtractor_0/XOR_3/NAND_2/a_6_n14# Gnd 0.14fF
C2202 addersubtractor_0/XOR_3/NAND_2/w_32_0# Gnd 0.40fF
C2203 addersubtractor_0/XOR_3/NAND_2/w_0_0# Gnd 0.40fF
C2204 addersubtractor_0/XOR_3/NAND_1/a_6_n14# Gnd 0.14fF
C2205 addersubtractor_0/XOR_3/NAND_3/in1 Gnd 0.78fF
C2206 addersubtractor_0/XOR_3/NAND_1/w_32_0# Gnd 0.40fF
C2207 addersubtractor_0/XOR_3/NAND_1/w_0_0# Gnd 0.40fF
C2208 addersubtractor_0/XOR_3/NAND_0/a_6_n14# Gnd 0.14fF
C2209 addersubtractor_0/XOR_3/NAND_2/in1 Gnd 0.97fF
C2210 addersubtractor_0/XOR_3/NAND_0/w_32_0# Gnd 0.40fF
C2211 addersubtractor_0/XOR_3/NAND_0/w_0_0# Gnd 0.40fF
C2212 addersubtractor_0/XOR_2/NAND_3/a_6_n14# Gnd 0.14fF
C2213 addersubtractor_0/XOR_2/NAND_3/in2 Gnd 0.76fF
C2214 addersubtractor_0/XOR_2/NAND_3/w_32_0# Gnd 0.40fF
C2215 addersubtractor_0/XOR_2/NAND_3/w_0_0# Gnd 0.40fF
C2216 addersubtractor_0/XOR_2/NAND_2/a_6_n14# Gnd 0.14fF
C2217 addersubtractor_0/XOR_2/NAND_2/w_32_0# Gnd 0.40fF
C2218 addersubtractor_0/XOR_2/NAND_2/w_0_0# Gnd 0.40fF
C2219 addersubtractor_0/XOR_2/NAND_1/a_6_n14# Gnd 0.14fF
C2220 addersubtractor_0/XOR_2/NAND_3/in1 Gnd 0.78fF
C2221 addersubtractor_0/XOR_2/NAND_1/w_32_0# Gnd 0.40fF
C2222 addersubtractor_0/XOR_2/NAND_1/w_0_0# Gnd 0.40fF
C2223 addersubtractor_0/XOR_2/NAND_0/a_6_n14# Gnd 0.14fF
C2224 addersubtractor_0/XOR_2/NAND_2/in1 Gnd 0.97fF
C2225 addersubtractor_0/XOR_2/NAND_0/w_32_0# Gnd 0.40fF
C2226 addersubtractor_0/XOR_2/NAND_0/w_0_0# Gnd 0.40fF
C2227 addersubtractor_0/XOR_1/NAND_3/a_6_n14# Gnd 0.14fF
C2228 addersubtractor_0/XOR_1/NAND_3/in2 Gnd 0.76fF
C2229 addersubtractor_0/XOR_1/NAND_3/w_32_0# Gnd 0.40fF
C2230 addersubtractor_0/XOR_1/NAND_3/w_0_0# Gnd 0.40fF
C2231 addersubtractor_0/XOR_1/NAND_2/a_6_n14# Gnd 0.14fF
C2232 addersubtractor_0/XOR_1/NAND_2/w_32_0# Gnd 0.40fF
C2233 addersubtractor_0/XOR_1/NAND_2/w_0_0# Gnd 0.40fF
C2234 addersubtractor_0/XOR_1/NAND_1/a_6_n14# Gnd 0.14fF
C2235 addersubtractor_0/XOR_1/NAND_3/in1 Gnd 0.78fF
C2236 addersubtractor_0/XOR_1/NAND_1/w_32_0# Gnd 0.40fF
C2237 addersubtractor_0/XOR_1/NAND_1/w_0_0# Gnd 0.40fF
C2238 addersubtractor_0/XOR_1/NAND_0/a_6_n14# Gnd 0.14fF
C2239 addersubtractor_0/XOR_1/NAND_2/in1 Gnd 0.97fF
C2240 addersubtractor_0/XOR_1/NAND_0/w_32_0# Gnd 0.40fF
C2241 addersubtractor_0/XOR_1/NAND_0/w_0_0# Gnd 0.40fF
C2242 addersubtractor_0/XOR_0/NAND_3/a_6_n14# Gnd 0.14fF
C2243 addersubtractor_0/XOR_0/NAND_3/in2 Gnd 0.76fF
C2244 addersubtractor_0/XOR_0/NAND_3/w_32_0# Gnd 0.40fF
C2245 addersubtractor_0/XOR_0/NAND_3/w_0_0# Gnd 0.40fF
C2246 addersubtractor_0/XOR_0/NAND_2/a_6_n14# Gnd 0.14fF
C2247 addersubtractor_0/XOR_0/NAND_2/w_32_0# Gnd 0.40fF
C2248 addersubtractor_0/XOR_0/NAND_2/w_0_0# Gnd 0.40fF
C2249 addersubtractor_0/XOR_0/NAND_1/a_6_n14# Gnd 0.14fF
C2250 addersubtractor_0/XOR_0/NAND_3/in1 Gnd 0.78fF
C2251 addersubtractor_0/XOR_0/NAND_1/w_32_0# Gnd 0.40fF
C2252 addersubtractor_0/XOR_0/NAND_1/w_0_0# Gnd 0.40fF
C2253 addersubtractor_0/XOR_0/NAND_0/a_6_n14# Gnd 0.14fF
C2254 addersubtractor_0/XOR_0/NAND_2/in1 Gnd 0.97fF
C2255 S0 Gnd 10.27fF
C2256 addersubtractor_0/XOR_0/NAND_0/w_32_0# Gnd 0.40fF
C2257 addersubtractor_0/XOR_0/NAND_0/w_0_0# Gnd 0.40fF
C2258 addersubtractor_0/fulladder_3/XOR_1/NAND_3/a_6_n14# Gnd 0.14fF
C2259 adder3 Gnd 0.51fF
C2260 addersubtractor_0/fulladder_3/XOR_1/NAND_3/in2 Gnd 0.76fF
C2261 addersubtractor_0/fulladder_3/XOR_1/NAND_3/w_32_0# Gnd 0.40fF
C2262 addersubtractor_0/fulladder_3/XOR_1/NAND_3/w_0_0# Gnd 0.40fF
C2263 addersubtractor_0/fulladder_3/XOR_1/NAND_2/a_6_n14# Gnd 0.14fF
C2264 addersubtractor_0/fulladder_3/XOR_1/NAND_2/w_32_0# Gnd 0.40fF
C2265 addersubtractor_0/fulladder_3/XOR_1/NAND_2/w_0_0# Gnd 0.40fF
C2266 addersubtractor_0/fulladder_3/XOR_1/NAND_1/a_6_n14# Gnd 0.14fF
C2267 addersubtractor_0/fulladder_3/XOR_1/NAND_3/in1 Gnd 0.78fF
C2268 addersubtractor_0/fulladder_3/XOR_1/NAND_1/w_32_0# Gnd 0.40fF
C2269 addersubtractor_0/fulladder_3/XOR_1/NAND_1/w_0_0# Gnd 0.40fF
C2270 addersubtractor_0/fulladder_3/XOR_1/NAND_0/a_6_n14# Gnd 0.14fF
C2271 addersubtractor_0/fulladder_3/XOR_1/NAND_2/in1 Gnd 0.97fF
C2272 addersubtractor_0/fulladder_2/C Gnd 1.24fF
C2273 addersubtractor_0/fulladder_3/XOR_1/NAND_0/w_32_0# Gnd 0.40fF
C2274 addersubtractor_0/fulladder_3/XOR_1/NAND_0/w_0_0# Gnd 0.40fF
C2275 addersubtractor_0/fulladder_3/OR_0/NOR_0/a_13_6# Gnd 0.02fF
C2276 addersubtractor_0/fulladder_3/OR_0/in1 Gnd 0.40fF
C2277 addersubtractor_0/fulladder_3/OR_0/NOR_0/w_32_0# Gnd 0.40fF
C2278 addersubtractor_0/fulladder_3/OR_0/NOR_0/w_0_0# Gnd 0.40fF
C2279 AND_0/in1 Gnd 0.43fF
C2280 addersubtractor_0/fulladder_3/OR_0/NOT_0/in Gnd 0.77fF
C2281 addersubtractor_0/fulladder_3/OR_0/NOT_0/w_0_0# Gnd 0.40fF
C2282 addersubtractor_0/fulladder_3/XOR_0/NAND_3/a_6_n14# Gnd 0.14fF
C2283 addersubtractor_0/fulladder_3/XOR_1/in2 Gnd 2.44fF
C2284 addersubtractor_0/fulladder_3/XOR_0/NAND_3/in2 Gnd 0.76fF
C2285 addersubtractor_0/fulladder_3/XOR_0/NAND_3/w_32_0# Gnd 0.40fF
C2286 addersubtractor_0/fulladder_3/XOR_0/NAND_3/w_0_0# Gnd 0.40fF
C2287 addersubtractor_0/fulladder_3/XOR_0/NAND_2/a_6_n14# Gnd 0.14fF
C2288 addersubtractor_0/fulladder_3/XOR_0/NAND_2/w_32_0# Gnd 0.40fF
C2289 addersubtractor_0/fulladder_3/XOR_0/NAND_2/w_0_0# Gnd 0.40fF
C2290 addersubtractor_0/fulladder_3/XOR_0/NAND_1/a_6_n14# Gnd 0.14fF
C2291 addersubtractor_0/fulladder_3/XOR_0/NAND_3/in1 Gnd 0.78fF
C2292 addersubtractor_0/fulladder_3/XOR_0/NAND_1/w_32_0# Gnd 0.40fF
C2293 addersubtractor_0/fulladder_3/XOR_0/NAND_1/w_0_0# Gnd 0.40fF
C2294 addersubtractor_0/fulladder_3/XOR_0/NAND_0/a_6_n14# Gnd 0.14fF
C2295 addersubtractor_0/fulladder_3/XOR_0/NAND_2/in1 Gnd 0.97fF
C2296 addersubtractor_0/XOR_3/out Gnd 1.88fF
C2297 enableblock_0/B_out1 Gnd 2.66fF
C2298 addersubtractor_0/fulladder_3/XOR_0/NAND_0/w_32_0# Gnd 0.40fF
C2299 addersubtractor_0/fulladder_3/XOR_0/NAND_0/w_0_0# Gnd 0.40fF
C2300 addersubtractor_0/fulladder_3/AND_1/not_0/in Gnd 0.76fF
C2301 addersubtractor_0/fulladder_3/AND_1/not_0/w_0_0# Gnd 0.40fF
C2302 addersubtractor_0/fulladder_3/AND_1/NAND_0/a_6_n14# Gnd 0.14fF
C2303 addersubtractor_0/fulladder_3/AND_1/NAND_0/w_32_0# Gnd 0.40fF
C2304 addersubtractor_0/fulladder_3/AND_1/NAND_0/w_0_0# Gnd 0.40fF
C2305 addersubtractor_0/fulladder_3/AND_0/not_0/in Gnd 0.76fF
C2306 addersubtractor_0/fulladder_3/OR_0/in2 Gnd 0.47fF
C2307 addersubtractor_0/fulladder_3/AND_0/not_0/w_0_0# Gnd 0.40fF
C2308 addersubtractor_0/fulladder_3/AND_0/NAND_0/a_6_n14# Gnd 0.14fF
C2309 addersubtractor_0/fulladder_3/AND_0/NAND_0/w_32_0# Gnd 0.40fF
C2310 addersubtractor_0/fulladder_3/AND_0/NAND_0/w_0_0# Gnd 0.40fF
C2311 addersubtractor_0/fulladder_2/XOR_1/NAND_3/a_6_n14# Gnd 0.14fF
C2312 adder2 Gnd 0.57fF
C2313 addersubtractor_0/fulladder_2/XOR_1/NAND_3/in2 Gnd 0.76fF
C2314 addersubtractor_0/fulladder_2/XOR_1/NAND_3/w_32_0# Gnd 0.40fF
C2315 addersubtractor_0/fulladder_2/XOR_1/NAND_3/w_0_0# Gnd 0.40fF
C2316 addersubtractor_0/fulladder_2/XOR_1/NAND_2/a_6_n14# Gnd 0.14fF
C2317 addersubtractor_0/fulladder_2/XOR_1/NAND_2/w_32_0# Gnd 0.40fF
C2318 addersubtractor_0/fulladder_2/XOR_1/NAND_2/w_0_0# Gnd 0.40fF
C2319 addersubtractor_0/fulladder_2/XOR_1/NAND_1/a_6_n14# Gnd 0.14fF
C2320 addersubtractor_0/fulladder_2/XOR_1/NAND_3/in1 Gnd 0.78fF
C2321 addersubtractor_0/fulladder_2/XOR_1/NAND_1/w_32_0# Gnd 0.40fF
C2322 addersubtractor_0/fulladder_2/XOR_1/NAND_1/w_0_0# Gnd 0.40fF
C2323 gnd Gnd 93.17fF
C2324 addersubtractor_0/fulladder_2/XOR_1/NAND_0/a_6_n14# Gnd 0.14fF
C2325 addersubtractor_0/fulladder_2/XOR_1/NAND_2/in1 Gnd 0.97fF
C2326 addersubtractor_0/fulladder_1/C Gnd 1.25fF
C2327 addersubtractor_0/fulladder_2/XOR_1/NAND_0/w_32_0# Gnd 0.40fF
C2328 addersubtractor_0/fulladder_2/XOR_1/NAND_0/w_0_0# Gnd 0.40fF
C2329 addersubtractor_0/fulladder_2/OR_0/NOR_0/a_13_6# Gnd 0.02fF
C2330 addersubtractor_0/fulladder_2/OR_0/in1 Gnd 0.40fF
C2331 addersubtractor_0/fulladder_2/OR_0/NOR_0/w_32_0# Gnd 0.40fF
C2332 addersubtractor_0/fulladder_2/OR_0/NOR_0/w_0_0# Gnd 0.40fF
C2333 addersubtractor_0/fulladder_2/OR_0/NOT_0/in Gnd 0.77fF
C2334 addersubtractor_0/fulladder_2/OR_0/NOT_0/w_0_0# Gnd 0.40fF
C2335 addersubtractor_0/fulladder_2/XOR_0/NAND_3/a_6_n14# Gnd 0.14fF
C2336 addersubtractor_0/fulladder_2/XOR_1/in2 Gnd 2.44fF
C2337 addersubtractor_0/fulladder_2/XOR_0/NAND_3/in2 Gnd 0.76fF
C2338 addersubtractor_0/fulladder_2/XOR_0/NAND_3/w_32_0# Gnd 0.40fF
C2339 addersubtractor_0/fulladder_2/XOR_0/NAND_3/w_0_0# Gnd 0.40fF
C2340 addersubtractor_0/fulladder_2/XOR_0/NAND_2/a_6_n14# Gnd 0.14fF
C2341 addersubtractor_0/fulladder_2/XOR_0/NAND_2/w_32_0# Gnd 0.40fF
C2342 addersubtractor_0/fulladder_2/XOR_0/NAND_2/w_0_0# Gnd 0.40fF
C2343 addersubtractor_0/fulladder_2/XOR_0/NAND_1/a_6_n14# Gnd 0.14fF
C2344 addersubtractor_0/fulladder_2/XOR_0/NAND_3/in1 Gnd 0.78fF
C2345 addersubtractor_0/fulladder_2/XOR_0/NAND_1/w_32_0# Gnd 0.40fF
C2346 addersubtractor_0/fulladder_2/XOR_0/NAND_1/w_0_0# Gnd 0.40fF
C2347 addersubtractor_0/fulladder_2/XOR_0/NAND_0/a_6_n14# Gnd 0.14fF
C2348 addersubtractor_0/fulladder_2/XOR_0/NAND_2/in1 Gnd 0.97fF
C2349 addersubtractor_0/XOR_2/out Gnd 1.88fF
C2350 enableblock_0/B_out3 Gnd 2.50fF
C2351 addersubtractor_0/fulladder_2/XOR_0/NAND_0/w_32_0# Gnd 0.40fF
C2352 addersubtractor_0/fulladder_2/XOR_0/NAND_0/w_0_0# Gnd 0.40fF
C2353 addersubtractor_0/fulladder_2/AND_1/not_0/in Gnd 0.76fF
C2354 addersubtractor_0/fulladder_2/AND_1/not_0/w_0_0# Gnd 0.40fF
C2355 addersubtractor_0/fulladder_2/AND_1/NAND_0/a_6_n14# Gnd 0.14fF
C2356 addersubtractor_0/fulladder_2/AND_1/NAND_0/w_32_0# Gnd 0.40fF
C2357 addersubtractor_0/fulladder_2/AND_1/NAND_0/w_0_0# Gnd 0.40fF
C2358 addersubtractor_0/fulladder_2/AND_0/not_0/in Gnd 0.76fF
C2359 addersubtractor_0/fulladder_2/OR_0/in2 Gnd 0.47fF
C2360 addersubtractor_0/fulladder_2/AND_0/not_0/w_0_0# Gnd 0.40fF
C2361 addersubtractor_0/fulladder_2/AND_0/NAND_0/a_6_n14# Gnd 0.14fF
C2362 addersubtractor_0/fulladder_2/AND_0/NAND_0/w_32_0# Gnd 0.40fF
C2363 addersubtractor_0/fulladder_2/AND_0/NAND_0/w_0_0# Gnd 0.40fF
C2364 addersubtractor_0/fulladder_1/XOR_1/NAND_3/a_6_n14# Gnd 0.14fF
C2365 adder1 Gnd 0.54fF
C2366 addersubtractor_0/fulladder_1/XOR_1/NAND_3/in2 Gnd 0.76fF
C2367 addersubtractor_0/fulladder_1/XOR_1/NAND_3/w_32_0# Gnd 0.40fF
C2368 addersubtractor_0/fulladder_1/XOR_1/NAND_3/w_0_0# Gnd 0.40fF
C2369 addersubtractor_0/fulladder_1/XOR_1/NAND_2/a_6_n14# Gnd 0.14fF
C2370 addersubtractor_0/fulladder_1/XOR_1/NAND_2/w_32_0# Gnd 0.40fF
C2371 addersubtractor_0/fulladder_1/XOR_1/NAND_2/w_0_0# Gnd 0.40fF
C2372 addersubtractor_0/fulladder_1/XOR_1/NAND_1/a_6_n14# Gnd 0.14fF
C2373 addersubtractor_0/fulladder_1/XOR_1/NAND_3/in1 Gnd 0.78fF
C2374 addersubtractor_0/fulladder_1/XOR_1/NAND_1/w_32_0# Gnd 0.40fF
C2375 addersubtractor_0/fulladder_1/XOR_1/NAND_1/w_0_0# Gnd 0.40fF
C2376 addersubtractor_0/fulladder_1/XOR_1/NAND_0/a_6_n14# Gnd 0.14fF
C2377 addersubtractor_0/fulladder_1/XOR_1/NAND_2/in1 Gnd 0.97fF
C2378 addersubtractor_0/fulladder_0/C Gnd 1.23fF
C2379 addersubtractor_0/fulladder_1/XOR_1/NAND_0/w_32_0# Gnd 0.40fF
C2380 addersubtractor_0/fulladder_1/XOR_1/NAND_0/w_0_0# Gnd 0.40fF
C2381 addersubtractor_0/fulladder_1/OR_0/NOR_0/a_13_6# Gnd 0.02fF
C2382 addersubtractor_0/fulladder_1/OR_0/in1 Gnd 0.40fF
C2383 addersubtractor_0/fulladder_1/OR_0/NOR_0/w_32_0# Gnd 0.40fF
C2384 addersubtractor_0/fulladder_1/OR_0/NOR_0/w_0_0# Gnd 0.40fF
C2385 addersubtractor_0/fulladder_1/OR_0/NOT_0/in Gnd 0.77fF
C2386 addersubtractor_0/fulladder_1/OR_0/NOT_0/w_0_0# Gnd 0.40fF
C2387 addersubtractor_0/fulladder_1/XOR_0/NAND_3/a_6_n14# Gnd 0.14fF
C2388 addersubtractor_0/fulladder_1/XOR_1/in2 Gnd 2.44fF
C2389 addersubtractor_0/fulladder_1/XOR_0/NAND_3/in2 Gnd 0.76fF
C2390 addersubtractor_0/fulladder_1/XOR_0/NAND_3/w_32_0# Gnd 0.40fF
C2391 addersubtractor_0/fulladder_1/XOR_0/NAND_3/w_0_0# Gnd 0.40fF
C2392 addersubtractor_0/fulladder_1/XOR_0/NAND_2/a_6_n14# Gnd 0.14fF
C2393 addersubtractor_0/fulladder_1/XOR_0/NAND_2/w_32_0# Gnd 0.40fF
C2394 addersubtractor_0/fulladder_1/XOR_0/NAND_2/w_0_0# Gnd 0.40fF
C2395 addersubtractor_0/fulladder_1/XOR_0/NAND_1/a_6_n14# Gnd 0.14fF
C2396 addersubtractor_0/fulladder_1/XOR_0/NAND_3/in1 Gnd 0.78fF
C2397 addersubtractor_0/fulladder_1/XOR_0/NAND_1/w_32_0# Gnd 0.40fF
C2398 addersubtractor_0/fulladder_1/XOR_0/NAND_1/w_0_0# Gnd 0.40fF
C2399 addersubtractor_0/fulladder_1/XOR_0/NAND_0/a_6_n14# Gnd 0.14fF
C2400 addersubtractor_0/fulladder_1/XOR_0/NAND_2/in1 Gnd 0.97fF
C2401 addersubtractor_0/XOR_1/out Gnd 1.88fF
C2402 enableblock_0/A_out1 Gnd 2.48fF
C2403 addersubtractor_0/fulladder_1/XOR_0/NAND_0/w_32_0# Gnd 0.40fF
C2404 addersubtractor_0/fulladder_1/XOR_0/NAND_0/w_0_0# Gnd 0.40fF
C2405 addersubtractor_0/fulladder_1/AND_1/not_0/in Gnd 0.76fF
C2406 addersubtractor_0/fulladder_1/AND_1/not_0/w_0_0# Gnd 0.40fF
C2407 addersubtractor_0/fulladder_1/AND_1/NAND_0/a_6_n14# Gnd 0.14fF
C2408 addersubtractor_0/fulladder_1/AND_1/NAND_0/w_32_0# Gnd 0.40fF
C2409 addersubtractor_0/fulladder_1/AND_1/NAND_0/w_0_0# Gnd 0.40fF
C2410 addersubtractor_0/fulladder_1/AND_0/not_0/in Gnd 0.76fF
C2411 addersubtractor_0/fulladder_1/OR_0/in2 Gnd 0.47fF
C2412 addersubtractor_0/fulladder_1/AND_0/not_0/w_0_0# Gnd 0.40fF
C2413 addersubtractor_0/fulladder_1/AND_0/NAND_0/a_6_n14# Gnd 0.14fF
C2414 addersubtractor_0/fulladder_1/AND_0/NAND_0/w_32_0# Gnd 0.40fF
C2415 addersubtractor_0/fulladder_1/AND_0/NAND_0/w_0_0# Gnd 0.40fF
C2416 addersubtractor_0/fulladder_0/XOR_1/NAND_3/a_6_n14# Gnd 0.14fF
C2417 adder0 Gnd 0.57fF
C2418 addersubtractor_0/fulladder_0/XOR_1/NAND_3/in2 Gnd 0.76fF
C2419 addersubtractor_0/fulladder_0/XOR_1/NAND_3/w_32_0# Gnd 0.40fF
C2420 addersubtractor_0/fulladder_0/XOR_1/NAND_3/w_0_0# Gnd 0.40fF
C2421 addersubtractor_0/fulladder_0/XOR_1/NAND_2/a_6_n14# Gnd 0.14fF
C2422 addersubtractor_0/fulladder_0/XOR_1/NAND_2/w_32_0# Gnd 0.40fF
C2423 addersubtractor_0/fulladder_0/XOR_1/NAND_2/w_0_0# Gnd 0.40fF
C2424 addersubtractor_0/fulladder_0/XOR_1/NAND_1/a_6_n14# Gnd 0.14fF
C2425 addersubtractor_0/fulladder_0/XOR_1/NAND_3/in1 Gnd 0.78fF
C2426 addersubtractor_0/fulladder_0/XOR_1/NAND_1/w_32_0# Gnd 0.40fF
C2427 addersubtractor_0/fulladder_0/XOR_1/NAND_1/w_0_0# Gnd 0.40fF
C2428 addersubtractor_0/fulladder_0/XOR_1/NAND_0/a_6_n14# Gnd 0.14fF
C2429 addersubtractor_0/fulladder_0/XOR_1/NAND_2/in1 Gnd 0.97fF
C2430 addersubtractor_0/fulladder_0/XOR_1/NAND_0/w_32_0# Gnd 0.40fF
C2431 addersubtractor_0/fulladder_0/XOR_1/NAND_0/w_0_0# Gnd 0.40fF
C2432 addersubtractor_0/fulladder_0/OR_0/NOR_0/a_13_6# Gnd 0.02fF
C2433 addersubtractor_0/fulladder_0/OR_0/in1 Gnd 0.40fF
C2434 addersubtractor_0/fulladder_0/OR_0/NOR_0/w_32_0# Gnd 0.40fF
C2435 addersubtractor_0/fulladder_0/OR_0/NOR_0/w_0_0# Gnd 0.40fF
C2436 addersubtractor_0/fulladder_0/OR_0/NOT_0/in Gnd 0.77fF
C2437 addersubtractor_0/fulladder_0/OR_0/NOT_0/w_0_0# Gnd 0.40fF
C2438 vdd Gnd 28.56fF
C2439 addersubtractor_0/fulladder_0/XOR_0/NAND_3/a_6_n14# Gnd 0.14fF
C2440 addersubtractor_0/fulladder_0/XOR_1/in2 Gnd 2.44fF
C2441 addersubtractor_0/fulladder_0/XOR_0/NAND_3/in2 Gnd 0.76fF
C2442 addersubtractor_0/fulladder_0/XOR_0/NAND_3/w_32_0# Gnd 0.40fF
C2443 addersubtractor_0/fulladder_0/XOR_0/NAND_3/w_0_0# Gnd 0.40fF
C2444 addersubtractor_0/fulladder_0/XOR_0/NAND_2/a_6_n14# Gnd 0.14fF
C2445 addersubtractor_0/fulladder_0/XOR_0/NAND_2/w_32_0# Gnd 0.40fF
C2446 addersubtractor_0/fulladder_0/XOR_0/NAND_2/w_0_0# Gnd 0.40fF
C2447 addersubtractor_0/fulladder_0/XOR_0/NAND_1/a_6_n14# Gnd 0.14fF
C2448 addersubtractor_0/fulladder_0/XOR_0/NAND_3/in1 Gnd 0.78fF
C2449 addersubtractor_0/fulladder_0/XOR_0/NAND_1/w_32_0# Gnd 0.40fF
C2450 addersubtractor_0/fulladder_0/XOR_0/NAND_1/w_0_0# Gnd 0.40fF
C2451 addersubtractor_0/fulladder_0/XOR_0/NAND_0/a_6_n14# Gnd 0.14fF
C2452 addersubtractor_0/fulladder_0/XOR_0/NAND_2/in1 Gnd 0.97fF
C2453 addersubtractor_0/XOR_0/out Gnd 1.87fF
C2454 enableblock_0/A_out3 Gnd 3.35fF
C2455 addersubtractor_0/fulladder_0/XOR_0/NAND_0/w_32_0# Gnd 0.40fF
C2456 addersubtractor_0/fulladder_0/XOR_0/NAND_0/w_0_0# Gnd 0.40fF
C2457 addersubtractor_0/fulladder_0/AND_1/not_0/in Gnd 0.76fF
C2458 addersubtractor_0/fulladder_0/AND_1/not_0/w_0_0# Gnd 0.40fF
C2459 addersubtractor_0/fulladder_0/AND_1/NAND_0/a_6_n14# Gnd 0.14fF
C2460 addersubtractor_0/fulladder_0/AND_1/NAND_0/w_32_0# Gnd 0.40fF
C2461 addersubtractor_0/fulladder_0/AND_1/NAND_0/w_0_0# Gnd 0.40fF
C2462 addersubtractor_0/fulladder_0/AND_0/not_0/in Gnd 0.76fF
C2463 addersubtractor_0/fulladder_0/OR_0/in2 Gnd 0.47fF
C2464 addersubtractor_0/fulladder_0/AND_0/not_0/w_0_0# Gnd 0.40fF
C2465 addersubtractor_0/fulladder_0/AND_0/NAND_0/a_6_n14# Gnd 0.14fF
C2466 addersubtractor_0/fulladder_0/AND_0/NAND_0/w_32_0# Gnd 0.40fF
C2467 vdd Gnd 0.40fF



.tran 1n 400n
*target text
.control
run
*quit
set color0 = rgb:f/f/e
set color1 = black
plot v(A0) v(A1)+2 v(A2)+4 v(A3)+6 v(B0)+8 v(B1)+10 v(B2)+12 v(B3)+14
plot v(S0) v(S1)+2 v(adder0)+4 v(adder1)+6 v(adder2)+8 v(adder3)+10 v(carry)+12
plot v(S0) v(S1)+2 v(lesser)+4 v(equal)+6 v(greater)+8 
plot v(S0) v(S1)+2 v(and0)+4 v(and1)+6 v(and2)+8 v(and3)+10 
.end
.endc