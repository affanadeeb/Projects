magic
tech scmos
timestamp 1698566035
<< nwell >>
rect 0 0 25 16
<< ntransistor >>
rect 11 -14 13 -10
<< ptransistor >>
rect 11 6 13 10
<< ndiffusion >>
rect 10 -14 11 -10
rect 13 -14 14 -10
<< pdiffusion >>
rect 10 6 11 10
rect 13 6 14 10
<< ndcontact >>
rect 6 -14 10 -10
rect 14 -14 18 -10
<< pdcontact >>
rect 6 6 10 10
rect 14 6 18 10
<< polysilicon >>
rect 11 10 13 13
rect 11 -3 13 6
rect 7 -7 13 -3
rect 11 -10 13 -7
rect 11 -17 13 -14
<< polycontact >>
rect 3 -7 7 -3
<< metal1 >>
rect 0 16 25 19
rect 7 10 10 16
rect 14 -3 17 6
rect 1 -7 3 -3
rect 14 -6 22 -3
rect 14 -10 17 -6
rect 7 -18 10 -14
rect 1 -21 25 -18
<< labels >>
rlabel metal1 0 16 25 19 5 vdd
rlabel metal1 17 -6 22 -3 1 out
rlabel metal1 1 -7 3 -3 3 in
rlabel metal1 1 -21 25 -18 1 gnd
<< end >>
